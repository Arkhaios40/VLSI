magic
tech sky130A
timestamp 1670361013
<< nwell >>
rect -279 -713 279 713
<< mvpmos >>
rect -150 -600 150 600
<< mvpdiff >>
rect -179 594 -150 600
rect -179 -594 -173 594
rect -156 -594 -150 594
rect -179 -600 -150 -594
rect 150 594 179 600
rect 150 -594 156 594
rect 173 -594 179 594
rect 150 -600 179 -594
<< mvpdiffc >>
rect -173 -594 -156 594
rect 156 -594 173 594
<< mvnsubdiff >>
rect -246 674 246 680
rect -246 657 -192 674
rect 192 657 246 674
rect -246 651 246 657
rect -246 626 -217 651
rect -246 -626 -240 626
rect -223 -626 -217 626
rect 217 626 246 651
rect -246 -651 -217 -626
rect 217 -626 223 626
rect 240 -626 246 626
rect 217 -651 246 -626
rect -246 -657 246 -651
rect -246 -674 -192 -657
rect 192 -674 246 -657
rect -246 -680 246 -674
<< mvnsubdiffcont >>
rect -192 657 192 674
rect -240 -626 -223 626
rect 223 -626 240 626
rect -192 -674 192 -657
<< poly >>
rect -150 600 150 613
rect -150 -613 150 -600
<< locali >>
rect -240 657 -192 674
rect 192 657 240 674
rect -240 626 -223 657
rect 223 626 240 657
rect -173 594 -156 602
rect -173 -602 -156 -594
rect 156 594 173 602
rect 156 -602 173 -594
rect -240 -657 -223 -626
rect 223 -657 240 -626
rect -240 -674 -192 -657
rect 192 -674 240 -657
<< viali >>
rect -173 -594 -156 594
rect 156 -594 173 594
<< metal1 >>
rect -176 594 -153 600
rect -176 -594 -173 594
rect -156 -594 -153 594
rect -176 -600 -153 -594
rect 153 594 176 600
rect 153 -594 156 594
rect 173 -594 176 594
rect 153 -600 176 -594
<< properties >>
string FIXED_BBOX -231 -665 231 665
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 12 l 3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
