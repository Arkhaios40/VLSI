magic
tech sky130A
magscale 1 2
timestamp 1669438545
<< pwell >>
rect -278 -2727 278 2727
<< mvnmos >>
rect -50 -2531 50 2469
<< mvndiff >>
rect -108 2457 -50 2469
rect -108 -2519 -96 2457
rect -62 -2519 -50 2457
rect -108 -2531 -50 -2519
rect 50 2457 108 2469
rect 50 -2519 62 2457
rect 96 -2519 108 2457
rect 50 -2531 108 -2519
<< mvndiffc >>
rect -96 -2519 -62 2457
rect 62 -2519 96 2457
<< mvpsubdiff >>
rect -242 2633 242 2691
rect -242 2583 -184 2633
rect -242 -2583 -230 2583
rect -196 -2583 -184 2583
rect 184 2583 242 2633
rect -242 -2633 -184 -2583
rect 184 -2583 196 2583
rect 230 -2583 242 2583
rect 184 -2633 242 -2583
rect -242 -2691 242 -2633
<< mvpsubdiffcont >>
rect -230 -2583 -196 2583
rect 196 -2583 230 2583
<< poly >>
rect -50 2541 50 2557
rect -50 2507 -34 2541
rect 34 2507 50 2541
rect -50 2469 50 2507
rect -50 -2557 50 -2531
<< polycont >>
rect -34 2507 34 2541
<< locali >>
rect -230 2583 -196 2607
rect 196 2583 230 2607
rect -50 2507 -34 2541
rect 34 2507 50 2541
rect -96 2457 -62 2473
rect -96 -2535 -62 -2519
rect 62 2457 96 2473
rect 62 -2535 96 -2519
rect -230 -2645 -196 -2583
rect 196 -2645 230 -2583
rect -230 -2679 230 -2645
<< viali >>
rect -34 2507 34 2541
rect -96 -2519 -62 2457
rect 62 -2519 96 2457
<< metal1 >>
rect -46 2541 46 2547
rect -46 2507 -34 2541
rect 34 2507 46 2541
rect -46 2501 46 2507
rect -102 2457 -56 2469
rect -102 -2519 -96 2457
rect -62 -2519 -56 2457
rect -102 -2531 -56 -2519
rect 56 2457 102 2469
rect 56 -2519 62 2457
rect 96 -2519 102 2457
rect 56 -2531 102 -2519
<< properties >>
string FIXED_BBOX -213 -2662 213 2662
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 25 l .5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
