magic
tech sky130A
timestamp 1669614457
<< mvnsubdiff >>
rect -1839 1918 -1810 2310
<< locali >>
rect -3912 3824 4052 3902
rect -3912 3385 -3805 3824
rect 3332 3385 4052 3824
rect -3912 3281 4052 3385
rect -506 2240 -242 3281
rect 3757 2269 4050 3281
rect -1736 2187 -242 2240
rect -1742 2064 -242 2187
rect -1736 2035 -242 2064
rect -1736 2029 -248 2035
rect 2673 2023 4050 2269
rect 2673 2017 4038 2023
rect 224 353 325 673
rect -4185 -22 -4089 300
rect 224 -22 329 353
rect -4185 -58 329 -22
rect -4185 -299 -3903 -58
rect -1490 -299 329 -58
rect -4185 -331 329 -299
rect -4185 -332 228 -331
rect -4185 -338 -4089 -332
<< viali >>
rect -3805 3385 3332 3824
rect -3903 -299 -1490 -58
<< metal1 >>
rect -1145 3901 915 3912
rect -1145 3892 3472 3901
rect -3891 3824 3472 3892
rect -3891 3385 -3805 3824
rect 3332 3385 3472 3824
rect -3891 3253 3472 3385
rect -3891 3110 -949 3253
rect 530 3119 3472 3253
rect -3915 -58 -1484 63
rect -3915 -299 -3903 -58
rect -1490 -299 -1484 -58
rect -3915 -631 -1484 -299
rect 507 -613 2920 45
use PMOSPair  PMOSPair_0
timestamp 1669589303
transform 1 0 424 0 1 -833
box -424 833 3216 4021
use PMOSPair  PMOSPair_1
timestamp 1669589303
transform 1 0 -3989 0 1 -830
box -424 833 3216 4021
<< labels >>
rlabel viali -3805 3385 3332 3824 1 Vss
port 0 n
rlabel metal1 515 -613 2898 -245 5 R_Pin
port 2 s
rlabel metal1 -3915 -631 -1484 -299 5 VP_LeftPin
port 1 s
<< end >>
