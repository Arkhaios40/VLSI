magic
tech sky130A
magscale 1 2
timestamp 1669447977
<< nwell >>
rect -758 -3262 758 3262
<< mvpmos >>
rect -500 -3036 500 2964
<< mvpdiff >>
rect -558 2952 -500 2964
rect -558 -3024 -546 2952
rect -512 -3024 -500 2952
rect -558 -3036 -500 -3024
rect 500 2952 558 2964
rect 500 -3024 512 2952
rect 546 -3024 558 2952
rect 500 -3036 558 -3024
<< mvpdiffc >>
rect -546 -3024 -512 2952
rect 512 -3024 546 2952
<< mvnsubdiff >>
rect -692 3138 692 3196
rect -692 3088 -634 3138
rect -692 -3088 -680 3088
rect -646 -3088 -634 3088
rect 634 3088 692 3138
rect -692 -3138 -634 -3088
rect 634 -3088 646 3088
rect 680 -3088 692 3088
rect 634 -3138 692 -3088
rect -692 -3196 692 -3138
<< mvnsubdiffcont >>
rect -680 -3088 -646 3088
rect 646 -3088 680 3088
<< poly >>
rect -500 3045 500 3061
rect -500 3011 -484 3045
rect 484 3011 500 3045
rect -500 2964 500 3011
rect -500 -3062 500 -3036
<< polycont >>
rect -484 3011 484 3045
<< locali >>
rect -398 3150 442 3184
rect 582 3150 680 3184
rect -680 3088 -646 3122
rect 646 3088 680 3150
rect -500 3011 -484 3045
rect 484 3011 500 3045
rect -546 2952 -512 2968
rect -546 -3040 -512 -3024
rect 512 2952 546 2968
rect 512 -3040 546 -3024
rect -680 -3138 -646 -3088
rect 646 -3138 680 -3088
<< viali >>
rect -546 -3024 -512 2952
rect 512 -3024 546 2952
<< metal1 >>
rect -552 2952 -506 2964
rect -552 -3024 -546 2952
rect -512 -3024 -506 2952
rect -552 -3036 -506 -3024
rect 506 2952 552 2964
rect 506 -3024 512 2952
rect 546 -3024 552 2952
rect 506 -3036 552 -3024
<< properties >>
string FIXED_BBOX -663 -3167 663 3167
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 30 l 5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
