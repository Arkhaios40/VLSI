magic
tech sky130A
magscale 1 2
timestamp 1669236281
<< pwell >>
rect -3898 -4598 3898 4598
<< psubdiff >>
rect -3862 4528 -3766 4562
rect 3766 4528 3862 4562
rect -3862 4466 -3828 4528
rect 3828 4466 3862 4528
rect -3862 -4528 -3828 -4466
rect 3828 -4528 3862 -4466
rect -3862 -4562 3862 -4528
<< psubdiffcont >>
rect -3766 4528 3766 4562
rect -3862 -4466 -3828 4466
rect 3828 -4466 3862 4466
<< xpolycontact >>
rect -3732 4000 -3450 4432
rect -3732 -4432 -3450 -4000
rect -3354 4000 -3072 4432
rect -3354 -4432 -3072 -4000
rect -2976 4000 -2694 4432
rect -2976 -4432 -2694 -4000
rect -2598 4000 -2316 4432
rect -2598 -4432 -2316 -4000
rect -2220 4000 -1938 4432
rect -2220 -4432 -1938 -4000
rect -1842 4000 -1560 4432
rect -1842 -4432 -1560 -4000
rect -1464 4000 -1182 4432
rect -1464 -4432 -1182 -4000
rect -1086 4000 -804 4432
rect -1086 -4432 -804 -4000
rect -708 4000 -426 4432
rect -708 -4432 -426 -4000
rect -330 4000 -48 4432
rect -330 -4432 -48 -4000
rect 48 4000 330 4432
rect 48 -4432 330 -4000
rect 426 4000 708 4432
rect 426 -4432 708 -4000
rect 804 4000 1086 4432
rect 804 -4432 1086 -4000
rect 1182 4000 1464 4432
rect 1182 -4432 1464 -4000
rect 1560 4000 1842 4432
rect 1560 -4432 1842 -4000
rect 1938 4000 2220 4432
rect 1938 -4432 2220 -4000
rect 2316 4000 2598 4432
rect 2316 -4432 2598 -4000
rect 2694 4000 2976 4432
rect 2694 -4432 2976 -4000
rect 3072 4000 3354 4432
rect 3072 -4432 3354 -4000
rect 3450 4000 3732 4432
rect 3450 -4432 3732 -4000
<< xpolyres >>
rect -3732 -4000 -3450 4000
rect -3354 -4000 -3072 4000
rect -2976 -4000 -2694 4000
rect -2598 -4000 -2316 4000
rect -2220 -4000 -1938 4000
rect -1842 -4000 -1560 4000
rect -1464 -4000 -1182 4000
rect -1086 -4000 -804 4000
rect -708 -4000 -426 4000
rect -330 -4000 -48 4000
rect 48 -4000 330 4000
rect 426 -4000 708 4000
rect 804 -4000 1086 4000
rect 1182 -4000 1464 4000
rect 1560 -4000 1842 4000
rect 1938 -4000 2220 4000
rect 2316 -4000 2598 4000
rect 2694 -4000 2976 4000
rect 3072 -4000 3354 4000
rect 3450 -4000 3732 4000
<< locali >>
rect -3862 4528 -3766 4562
rect 3766 4528 3862 4562
rect -3862 4466 -3828 4528
rect 3828 4466 3862 4528
rect -3862 -4528 -3828 -4466
rect 3828 -4528 3862 -4466
rect -3862 -4562 3862 -4528
<< viali >>
rect -3716 4017 -3466 4414
rect -3338 4017 -3088 4414
rect -2960 4017 -2710 4414
rect -2582 4017 -2332 4414
rect -2204 4017 -1954 4414
rect -1826 4017 -1576 4414
rect -1448 4017 -1198 4414
rect -1070 4017 -820 4414
rect -692 4017 -442 4414
rect -314 4017 -64 4414
rect 64 4017 314 4414
rect 442 4017 692 4414
rect 820 4017 1070 4414
rect 1198 4017 1448 4414
rect 1576 4017 1826 4414
rect 1954 4017 2204 4414
rect 2332 4017 2582 4414
rect 2710 4017 2960 4414
rect 3088 4017 3338 4414
rect 3466 4017 3716 4414
rect -3716 -4414 -3466 -4017
rect -3338 -4414 -3088 -4017
rect -2960 -4414 -2710 -4017
rect -2582 -4414 -2332 -4017
rect -2204 -4414 -1954 -4017
rect -1826 -4414 -1576 -4017
rect -1448 -4414 -1198 -4017
rect -1070 -4414 -820 -4017
rect -692 -4414 -442 -4017
rect -314 -4414 -64 -4017
rect 64 -4414 314 -4017
rect 442 -4414 692 -4017
rect 820 -4414 1070 -4017
rect 1198 -4414 1448 -4017
rect 1576 -4414 1826 -4017
rect 1954 -4414 2204 -4017
rect 2332 -4414 2582 -4017
rect 2710 -4414 2960 -4017
rect 3088 -4414 3338 -4017
rect 3466 -4414 3716 -4017
<< metal1 >>
rect -3722 4414 -3460 4426
rect -3722 4017 -3716 4414
rect -3466 4017 -3460 4414
rect -3722 4005 -3460 4017
rect -3344 4414 -3082 4426
rect -3344 4017 -3338 4414
rect -3088 4017 -3082 4414
rect -3344 4005 -3082 4017
rect -2966 4414 -2704 4426
rect -2966 4017 -2960 4414
rect -2710 4017 -2704 4414
rect -2966 4005 -2704 4017
rect -2588 4414 -2326 4426
rect -2588 4017 -2582 4414
rect -2332 4017 -2326 4414
rect -2588 4005 -2326 4017
rect -2210 4414 -1948 4426
rect -2210 4017 -2204 4414
rect -1954 4017 -1948 4414
rect -2210 4005 -1948 4017
rect -1832 4414 -1570 4426
rect -1832 4017 -1826 4414
rect -1576 4017 -1570 4414
rect -1832 4005 -1570 4017
rect -1454 4414 -1192 4426
rect -1454 4017 -1448 4414
rect -1198 4017 -1192 4414
rect -1454 4005 -1192 4017
rect -1076 4414 -814 4426
rect -1076 4017 -1070 4414
rect -820 4017 -814 4414
rect -1076 4005 -814 4017
rect -698 4414 -436 4426
rect -698 4017 -692 4414
rect -442 4017 -436 4414
rect -698 4005 -436 4017
rect -320 4414 -58 4426
rect -320 4017 -314 4414
rect -64 4017 -58 4414
rect -320 4005 -58 4017
rect 58 4414 320 4426
rect 58 4017 64 4414
rect 314 4017 320 4414
rect 58 4005 320 4017
rect 436 4414 698 4426
rect 436 4017 442 4414
rect 692 4017 698 4414
rect 436 4005 698 4017
rect 814 4414 1076 4426
rect 814 4017 820 4414
rect 1070 4017 1076 4414
rect 814 4005 1076 4017
rect 1192 4414 1454 4426
rect 1192 4017 1198 4414
rect 1448 4017 1454 4414
rect 1192 4005 1454 4017
rect 1570 4414 1832 4426
rect 1570 4017 1576 4414
rect 1826 4017 1832 4414
rect 1570 4005 1832 4017
rect 1948 4414 2210 4426
rect 1948 4017 1954 4414
rect 2204 4017 2210 4414
rect 1948 4005 2210 4017
rect 2326 4414 2588 4426
rect 2326 4017 2332 4414
rect 2582 4017 2588 4414
rect 2326 4005 2588 4017
rect 2704 4414 2966 4426
rect 2704 4017 2710 4414
rect 2960 4017 2966 4414
rect 2704 4005 2966 4017
rect 3082 4414 3344 4426
rect 3082 4017 3088 4414
rect 3338 4017 3344 4414
rect 3082 4005 3344 4017
rect 3460 4414 3722 4426
rect 3460 4017 3466 4414
rect 3716 4017 3722 4414
rect 3460 4005 3722 4017
rect -3722 -4017 -3460 -4005
rect -3722 -4414 -3716 -4017
rect -3466 -4414 -3460 -4017
rect -3722 -4426 -3460 -4414
rect -3344 -4017 -3082 -4005
rect -3344 -4414 -3338 -4017
rect -3088 -4414 -3082 -4017
rect -3344 -4426 -3082 -4414
rect -2966 -4017 -2704 -4005
rect -2966 -4414 -2960 -4017
rect -2710 -4414 -2704 -4017
rect -2966 -4426 -2704 -4414
rect -2588 -4017 -2326 -4005
rect -2588 -4414 -2582 -4017
rect -2332 -4414 -2326 -4017
rect -2588 -4426 -2326 -4414
rect -2210 -4017 -1948 -4005
rect -2210 -4414 -2204 -4017
rect -1954 -4414 -1948 -4017
rect -2210 -4426 -1948 -4414
rect -1832 -4017 -1570 -4005
rect -1832 -4414 -1826 -4017
rect -1576 -4414 -1570 -4017
rect -1832 -4426 -1570 -4414
rect -1454 -4017 -1192 -4005
rect -1454 -4414 -1448 -4017
rect -1198 -4414 -1192 -4017
rect -1454 -4426 -1192 -4414
rect -1076 -4017 -814 -4005
rect -1076 -4414 -1070 -4017
rect -820 -4414 -814 -4017
rect -1076 -4426 -814 -4414
rect -698 -4017 -436 -4005
rect -698 -4414 -692 -4017
rect -442 -4414 -436 -4017
rect -698 -4426 -436 -4414
rect -320 -4017 -58 -4005
rect -320 -4414 -314 -4017
rect -64 -4414 -58 -4017
rect -320 -4426 -58 -4414
rect 58 -4017 320 -4005
rect 58 -4414 64 -4017
rect 314 -4414 320 -4017
rect 58 -4426 320 -4414
rect 436 -4017 698 -4005
rect 436 -4414 442 -4017
rect 692 -4414 698 -4017
rect 436 -4426 698 -4414
rect 814 -4017 1076 -4005
rect 814 -4414 820 -4017
rect 1070 -4414 1076 -4017
rect 814 -4426 1076 -4414
rect 1192 -4017 1454 -4005
rect 1192 -4414 1198 -4017
rect 1448 -4414 1454 -4017
rect 1192 -4426 1454 -4414
rect 1570 -4017 1832 -4005
rect 1570 -4414 1576 -4017
rect 1826 -4414 1832 -4017
rect 1570 -4426 1832 -4414
rect 1948 -4017 2210 -4005
rect 1948 -4414 1954 -4017
rect 2204 -4414 2210 -4017
rect 1948 -4426 2210 -4414
rect 2326 -4017 2588 -4005
rect 2326 -4414 2332 -4017
rect 2582 -4414 2588 -4017
rect 2326 -4426 2588 -4414
rect 2704 -4017 2966 -4005
rect 2704 -4414 2710 -4017
rect 2960 -4414 2966 -4017
rect 2704 -4426 2966 -4414
rect 3082 -4017 3344 -4005
rect 3082 -4414 3088 -4017
rect 3338 -4414 3344 -4017
rect 3082 -4426 3344 -4414
rect 3460 -4017 3722 -4005
rect 3460 -4414 3466 -4017
rect 3716 -4414 3722 -4017
rect 3460 -4426 3722 -4414
<< res1p41 >>
rect -3734 -4002 -3448 4002
rect -3356 -4002 -3070 4002
rect -2978 -4002 -2692 4002
rect -2600 -4002 -2314 4002
rect -2222 -4002 -1936 4002
rect -1844 -4002 -1558 4002
rect -1466 -4002 -1180 4002
rect -1088 -4002 -802 4002
rect -710 -4002 -424 4002
rect -332 -4002 -46 4002
rect 46 -4002 332 4002
rect 424 -4002 710 4002
rect 802 -4002 1088 4002
rect 1180 -4002 1466 4002
rect 1558 -4002 1844 4002
rect 1936 -4002 2222 4002
rect 2314 -4002 2600 4002
rect 2692 -4002 2978 4002
rect 3070 -4002 3356 4002
rect 3448 -4002 3734 4002
<< properties >>
string FIXED_BBOX -3845 -4545 3845 4545
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 40 m 1 nx 20 wmin 1.410 lmin 0.50 rho 2000 val 57.004k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
