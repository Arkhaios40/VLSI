magic
tech sky130A
timestamp 1670432383
<< nwell >>
rect -1200 -90 3770 2650
<< locali >>
rect -770 2150 120 2190
rect -770 2070 -700 2150
rect 60 2070 120 2150
rect -770 2020 120 2070
rect 410 2100 2090 2310
rect 410 1940 500 2100
rect 410 1860 520 1940
rect 420 1573 510 1689
rect 420 1493 432 1573
rect 497 1493 510 1573
rect 420 1371 510 1493
rect 0 880 190 930
rect 410 890 510 1170
rect 1920 1093 2090 2100
rect 2330 2140 3310 2160
rect 2330 2030 2360 2140
rect 3280 2030 3310 2140
rect 2330 1990 3310 2030
rect 0 50 30 880
rect 170 838 190 880
rect 230 838 510 890
rect 170 560 510 838
rect 170 288 190 560
rect 230 288 510 560
rect 170 50 510 288
rect 0 20 510 50
rect 140 10 510 20
rect 230 -10 510 10
<< viali >>
rect -700 2070 60 2150
rect 432 1493 497 1573
rect 2360 2030 3280 2140
rect 30 50 170 880
<< metal1 >>
rect -800 2150 3390 2210
rect -800 2080 -700 2150
rect -799 2070 -700 2080
rect 60 2140 3390 2150
rect 60 2080 2360 2140
rect 60 2070 204 2080
rect -799 1953 204 2070
rect 704 1948 1707 2080
rect 2280 2030 2360 2080
rect 3280 2030 3390 2140
rect 2280 1930 3390 2030
rect -799 1580 204 1645
rect -799 1573 509 1580
rect -799 1493 432 1573
rect 497 1493 509 1573
rect -799 1476 509 1493
rect -799 1408 204 1476
rect 704 1397 1707 1637
rect 2320 1380 3323 1622
rect -800 880 200 1100
rect -800 509 30 880
rect -3826 182 30 509
rect -803 50 30 182
rect 170 50 200 880
rect 820 488 1520 1080
rect 2420 1069 3120 1080
rect 2217 742 4152 1069
rect 820 458 1521 488
rect 820 131 4151 458
rect 820 130 1515 131
rect 1362 122 1515 130
rect -803 28 200 50
rect -800 0 200 28
use sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ  sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_0
timestamp 1670432383
transform 0 1 -267 -1 0 1251
box -279 -731 279 856
use sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ  sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_1
timestamp 1670432383
transform 0 -1 1187 1 0 1242
box -279 -731 279 856
use sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ  sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_2
timestamp 1670432383
transform 0 1 -267 -1 0 1801
box -279 -731 279 856
use sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ  sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_3
timestamp 1670432383
transform 0 -1 2776 1 0 1229
box -279 -731 279 856
use sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ  sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_4
timestamp 1670432383
transform 0 -1 1194 1 0 1794
box -279 -731 279 856
use sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ  sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_5
timestamp 1670432383
transform 0 -1 2786 1 0 1769
box -279 -731 279 856
<< labels >>
rlabel metal1 -3826 182 30 509 7 In
port 0 w
rlabel metal1 2217 742 4152 1069 3 Cp1
port 1 e
rlabel metal1 820 131 4151 458 3 Cp2
port 2 e
<< end >>
