** sch_path: /home/arkhaios/Project/xschem/PrimalStructures/GainStage.sch
**.subckt GainStage Vplus Gain_L_Pin Gain_R_Pin Gate_Ref Out Gain_Vs
*.iopin Vplus
*.iopin Gain_L_Pin
*.iopin Gain_R_Pin
*.iopin Gate_Ref
*.iopin Out
*.iopin Gain_Vs
XM3 Out Gate_Ref Vplus Vplus sky130_fd_pr__pfet_g5v0d10v5 L=5 W=90 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Out Gain_R_Pin Gain_Vs Gain_Vs sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=50 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 Gain_R_Pin Gain_L_Pin Gain_Vs Gain_Vs sky130_fd_pr__nfet_g5v0d10v5 L=3 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 Gain_L_Pin Gain_L_Pin Gain_Vs Gain_Vs sky130_fd_pr__nfet_g5v0d10v5 L=3 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 Gain_R_Pin Out sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
**.ends
.end
