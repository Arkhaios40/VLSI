magic
tech sky130A
magscale 1 2
timestamp 1670983913
<< poly >>
rect 16200 26000 16800 26400
<< metal1 >>
rect -2468 52426 2938 53164
rect 4174 52316 11231 53054
rect 11969 52316 11975 53054
rect 13200 49234 15200 49400
rect 4560 47574 13370 49234
rect 15030 47574 15200 49234
rect 13200 47400 15200 47574
rect -2560 45618 2846 46356
rect 4008 45544 13431 46282
rect 14169 45544 14175 46282
rect 16400 42536 18400 42800
rect 4726 40876 16570 42536
rect 18230 40876 18400 42536
rect 16400 40600 18400 40876
rect -2654 38828 2752 39566
rect 3916 38828 15631 39566
rect 16369 38828 16375 39566
rect 19200 35728 21200 36000
rect 4580 34068 19370 35728
rect 21030 34068 21200 35728
rect 19200 33800 21200 34068
rect -2708 31964 2698 32702
rect 3620 32056 17831 32794
rect 18569 32056 18575 32794
rect 22000 28790 24000 29000
rect 4634 27130 22170 28790
rect 23830 27130 24000 28790
rect 22000 27000 24000 27130
rect -2728 25248 2678 25986
rect 3638 25230 8034 25968
rect 8769 25230 9044 25968
rect 4654 20360 6570 22020
rect 8230 20360 8326 22020
rect -2820 18404 2586 19142
rect 3472 18366 8031 19104
rect 8769 18366 8878 19104
rect 4726 13624 6738 15284
rect 8398 13624 8404 15284
rect -2948 11670 2458 12408
rect 3564 11632 8031 12370
rect 8769 11632 8970 12370
rect 6400 8642 8600 9000
rect 4672 6982 6684 8642
rect 8344 6982 8600 8642
rect 6400 6800 8600 6982
rect -3040 4860 2366 5598
rect 4008 4806 8431 5544
rect 9169 4806 9414 5544
rect 6600 1724 8600 2000
rect 4782 64 6794 1724
rect 8454 64 8600 1724
rect 6600 -200 8600 64
<< via1 >>
rect 11231 52316 11969 53054
rect 13370 47574 15030 49234
rect 13431 45544 14169 46282
rect 16570 40876 18230 42536
rect 15631 38828 16369 39566
rect 19370 34068 21030 35728
rect 17831 32056 18569 32794
rect 22170 27130 23830 28790
rect 8034 25230 8769 25968
rect 6570 20360 8230 22020
rect 8031 18366 8769 19104
rect 6738 13624 8398 15284
rect 8031 11632 8769 12370
rect 6684 6982 8344 8642
rect 8431 4806 9169 5544
rect 6794 64 8454 1724
<< metal2 >>
rect 20800 53167 22000 53400
rect 11232 53060 21032 53167
rect 11231 53054 21032 53060
rect 11969 52432 21032 53054
rect 21767 52432 22000 53167
rect 11231 52310 11969 52316
rect 8034 25968 8769 25974
rect 11232 25967 11967 52310
rect 20800 52200 22000 52432
rect 13200 49234 15200 49400
rect 13200 47574 13370 49234
rect 15030 47574 15200 49234
rect 13200 47400 15200 47574
rect 8769 25232 11967 25967
rect 13031 46282 21231 46369
rect 13031 45544 13431 46282
rect 14169 45631 21231 46282
rect 21969 45631 22369 46369
rect 13031 45538 14169 45544
rect 8034 25224 8769 25230
rect 6561 20360 6570 22020
rect 8230 20360 8239 22020
rect 8031 19104 8769 19110
rect 13031 19104 13769 45538
rect 16400 42536 18400 42800
rect 16400 40876 16570 42536
rect 18230 40876 18400 42536
rect 16400 40600 18400 40876
rect 15631 39569 16369 39572
rect 8769 18366 13769 19104
rect 15431 39566 21231 39569
rect 15431 38828 15631 39566
rect 16369 38831 21231 39566
rect 21969 38831 22369 39569
rect 15431 38822 16369 38828
rect 8031 18360 8769 18366
rect 6738 15284 8398 15290
rect 6729 13624 6738 15284
rect 8398 13624 8407 15284
rect 6738 13618 8398 13624
rect 8031 12370 8769 12376
rect 15431 12370 16169 38822
rect 19200 35728 21200 36000
rect 19200 34068 19370 35728
rect 21030 34068 21200 35728
rect 19200 33800 21200 34068
rect 8769 11632 16169 12370
rect 17831 32794 18569 32800
rect 24231 32769 24969 32778
rect 18569 32056 24231 32769
rect 17831 32031 24231 32056
rect 8031 11626 8769 11632
rect 6400 8642 8600 9000
rect 6400 6982 6684 8642
rect 8344 6982 8600 8642
rect 6400 6800 8600 6982
rect 8431 5544 9169 5550
rect 17831 5544 18569 32031
rect 24231 32022 24969 32031
rect 22000 28790 24000 29000
rect 22000 27130 22170 28790
rect 23830 27130 24000 28790
rect 22000 27000 24000 27130
rect 9169 4806 18569 5544
rect 8431 4800 9169 4806
rect 6600 1724 8600 2000
rect 6600 64 6794 1724
rect 8454 64 8600 1724
rect 6600 -200 8600 64
<< via2 >>
rect 21032 52432 21767 53167
rect 13370 47574 15030 49234
rect 21231 45631 21969 46369
rect 6570 20360 8230 22020
rect 16570 40876 18230 42536
rect 21231 38831 21969 39569
rect 6738 13624 8398 15284
rect 19370 34068 21030 35728
rect 24231 32031 24969 32769
rect 6684 6982 8344 8642
rect 22170 27130 23830 28790
rect 6794 64 8454 1724
<< metal3 >>
rect 21027 53167 21772 53172
rect 21027 52432 21032 53167
rect 21767 52432 28367 53167
rect 21027 52427 21772 52432
rect 13200 49234 15200 49400
rect 13200 47574 13370 49234
rect 15030 47574 15200 49234
rect 13200 47400 15200 47574
rect 13370 22030 15030 47400
rect 21226 46369 21974 46374
rect 21226 45631 21231 46369
rect 21969 45631 28369 46369
rect 21226 45626 21974 45631
rect 16400 42536 18400 42800
rect 16400 42531 16570 42536
rect 18230 42531 18400 42536
rect 16400 40871 16565 42531
rect 18235 40871 18400 42531
rect 16400 40600 18400 40871
rect 21226 39569 21974 39574
rect 21226 38831 21231 39569
rect 21969 38831 27769 39569
rect 21226 38826 21974 38831
rect 19200 35733 21200 36000
rect 19200 34063 19365 35733
rect 21035 34063 21200 35733
rect 19200 33800 21200 34063
rect 24226 32769 24974 32774
rect 24226 32031 24231 32769
rect 24969 32031 27769 32769
rect 24226 32026 24974 32031
rect 22000 28795 24000 29000
rect 22000 27125 22165 28795
rect 23835 27125 24000 28795
rect 22000 27000 24000 27125
rect 6565 22020 6575 22025
rect 6565 20360 6570 22020
rect 6565 20355 6575 20360
rect 8235 20355 8241 22025
rect 10970 20370 28030 22030
rect 6733 15284 8403 15289
rect 10970 15284 12630 20370
rect 6733 13624 6738 15284
rect 8398 13624 12630 15284
rect 13370 15229 28230 15230
rect 6733 13619 8403 13624
rect 13365 13571 13371 15229
rect 15029 15029 28230 15229
rect 15029 13571 16571 15029
rect 13370 13570 16571 13571
rect 16565 13371 16571 13570
rect 18229 13570 28230 15029
rect 18229 13371 18235 13570
rect 6400 8647 8600 9000
rect 6400 6977 6679 8647
rect 8349 6977 8600 8647
rect 19365 8630 19371 8829
rect 6400 6800 8600 6977
rect 11170 7171 19371 8630
rect 21029 8630 21035 8829
rect 21029 7171 28030 8630
rect 11170 6970 28030 7171
rect 6789 1724 8459 1729
rect 11170 1724 12830 6970
rect 22165 1830 22171 2029
rect 13570 1829 22171 1830
rect 6789 64 6794 1724
rect 8454 64 12830 1724
rect 13565 171 13571 1829
rect 15229 371 22171 1829
rect 23829 1830 23835 2029
rect 23829 371 27030 1830
rect 15229 171 27030 371
rect 13570 170 27030 171
rect 6789 59 8459 64
<< via3 >>
rect 16565 40876 16570 42531
rect 16570 40876 18230 42531
rect 18230 40876 18235 42531
rect 16565 40871 18235 40876
rect 19365 35728 21035 35733
rect 19365 34068 19370 35728
rect 19370 34068 21030 35728
rect 21030 34068 21035 35728
rect 19365 34063 21035 34068
rect 22165 28790 23835 28795
rect 22165 27130 22170 28790
rect 22170 27130 23830 28790
rect 23830 27130 23835 28790
rect 22165 27125 23835 27130
rect 6575 22020 8235 22025
rect 6575 20360 8230 22020
rect 8230 20360 8235 22020
rect 6575 20355 8235 20360
rect 13371 13571 15029 15229
rect 16571 13371 18229 15029
rect 6679 8642 8349 8647
rect 6679 6982 6684 8642
rect 6684 6982 8344 8642
rect 8344 6982 8349 8642
rect 6679 6977 8349 6982
rect 19371 7171 21029 8829
rect 13571 171 15229 1829
rect 22171 371 23829 2029
<< metal4 >>
rect 16564 42531 18236 42532
rect 16564 40871 16565 42531
rect 18235 40871 18236 42531
rect 16564 40870 18236 40871
rect 6574 22025 8236 22026
rect 6574 20355 6575 22025
rect 8235 22020 8236 22025
rect 8235 20360 10630 22020
rect 8235 20355 8236 20360
rect 6574 20354 8236 20355
rect 8970 17830 10630 20360
rect 8970 16170 15030 17830
rect 13370 15229 15030 16170
rect 13370 13571 13371 15229
rect 15029 13571 15030 15229
rect 13370 13570 15030 13571
rect 16570 15029 18230 40870
rect 19364 35733 21036 35734
rect 19364 34063 19365 35733
rect 21035 34063 21036 35733
rect 19364 34062 21036 34063
rect 16570 13371 16571 15029
rect 18229 13371 18230 15029
rect 16570 13370 18230 13371
rect 6400 8647 8600 9000
rect 6400 6977 6679 8647
rect 8349 8642 8600 8647
rect 19370 8829 21030 34062
rect 22164 28795 23836 28796
rect 22164 27125 22165 28795
rect 23835 27125 23836 28795
rect 22164 27124 23836 27125
rect 8349 6982 11630 8642
rect 19370 7171 19371 8829
rect 21029 7171 21030 8829
rect 19370 7170 21030 7171
rect 8349 6977 8600 6982
rect 6400 6800 8600 6977
rect 9970 4030 11630 6982
rect 9970 2370 15230 4030
rect 13570 1829 15230 2370
rect 13570 171 13571 1829
rect 15229 171 15230 1829
rect 22170 2029 23830 27124
rect 22170 371 22171 2029
rect 23829 371 23830 2029
rect 22170 370 23830 371
rect 13570 170 15230 171
use NmosStage1  NmosStage1_0
timestamp 1670981651
transform 1 0 4126 0 1 50852
box -3900 -3860 1854 2280
use NmosStage1  NmosStage1_1
timestamp 1670981651
transform 1 0 3830 0 1 3352
box -3900 -3860 1854 2280
use NmosStage1  NmosStage1_2
timestamp 1670981651
transform 1 0 3870 0 1 10198
box -3900 -3860 1854 2280
use NmosStage1  NmosStage1_3
timestamp 1670981651
transform 1 0 3852 0 1 16846
box -3900 -3860 1854 2280
use NmosStage1  NmosStage1_4
timestamp 1670981651
transform 1 0 3942 0 1 23676
box -3900 -3860 1854 2280
use NmosStage1  NmosStage1_5
timestamp 1670981651
transform 1 0 3942 0 1 30488
box -3900 -3860 1854 2280
use NmosStage1  NmosStage1_6
timestamp 1670981651
transform 1 0 3998 0 1 37302
box -3900 -3860 1854 2280
use NmosStage1  NmosStage1_7
timestamp 1670981651
transform 1 0 4034 0 1 44076
box -3900 -3860 1854 2280
<< labels >>
rlabel space 7000 52200 8400 53400 1 exists
rlabel metal1 -2200 52600 -1200 53000 7 Bit0i+
port 0 w
rlabel metal3 26600 52600 28000 53000 3 Out1
port 1 e
rlabel metal1 -2400 45800 -1000 46200 7 Bit0i-
port 2 w
rlabel metal3 26600 45800 28000 46200 3 Out2
port 3 e
rlabel metal1 -2400 39000 -1000 39400 7 Bit0q+
port 4 w
rlabel metal3 26200 39000 27600 39400 3 Out3
port 5 e
rlabel metal1 -2600 32200 -1200 32600 7 Bit0q-
port 6 w
rlabel metal3 26200 32200 27600 32600 3 Out4
port 7 e
rlabel metal1 -2600 25400 -1200 25800 7 Bit1i+
port 8 w
rlabel metal3 26200 21000 27600 21400 3 Out5
port 9 e
rlabel metal1 -2600 18600 -1200 19000 7 Bit1i-
port 10 w
rlabel metal3 26400 14200 27800 14600 3 Out6
port 11 e
rlabel metal1 -2600 11800 -1200 12200 7 bit1q+
port 12 w
rlabel metal3 26200 7600 27600 8000 3 Out7
port 13 e
rlabel metal1 -2600 5000 -1200 5400 7 Bit1q-
port 14 w
rlabel metal3 25200 800 26600 1200 3 Out8
port 15 e
<< end >>
