magic
tech sky130A
magscale 1 2
timestamp 1670907597
<< locali >>
rect -3780 260 -1180 500
rect -860 260 1740 500
rect -2120 -1200 -2000 -600
rect -2440 -1440 -2000 -1200
rect -2440 -3560 -2380 -1440
rect -2140 -2040 -2000 -1440
rect -2140 -3560 -2020 -2040
rect -2440 -3680 -2020 -3560
rect -1140 -3680 -880 -1140
rect -20 -2040 100 -600
<< viali >>
rect -2380 -3560 -2140 -1440
<< metal1 >>
rect -3700 1220 -1080 2280
rect -600 1220 1540 2280
rect -3700 1200 -780 1220
rect -1280 680 -780 1200
rect -3700 640 -780 680
rect -3700 120 -1060 640
rect -660 140 1560 620
rect -3700 60 -774 120
rect -1280 -460 -774 60
rect -1160 -820 -900 -460
rect -1860 -1040 -160 -820
rect -1860 -1220 -1300 -1040
rect -720 -1220 -160 -1040
rect -3660 -1440 -1854 -1340
rect -3660 -3560 -2380 -1440
rect -2140 -3560 -1854 -1440
rect -3660 -3680 -1854 -3560
rect -1260 -3620 -760 -1340
rect -140 -3660 1660 -1320
use sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z  sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_0
timestamp 1670907597
transform 0 -1 -2473 1 0 -172
box -528 -1427 528 1427
use sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z  sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_1
timestamp 1670907597
transform -1 0 -1572 0 -1 -2433
box -528 -1427 528 1427
use sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z  sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_2
timestamp 1670907597
transform 0 -1 -2473 1 0 928
box -528 -1427 528 1427
use sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z  sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_3
timestamp 1670907597
transform -1 0 -452 0 -1 -2433
box -528 -1427 528 1427
use sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z  sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_4
timestamp 1670907597
transform 0 1 427 -1 0 928
box -528 -1427 528 1427
use sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z  sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_5
timestamp 1670907597
transform 0 1 427 -1 0 -172
box -528 -1427 528 1427
<< labels >>
rlabel metal1 -3120 1700 -1760 2060 7 In
port 0 w
rlabel metal1 -220 1700 1120 2060 3 Cp1
port 1 e
rlabel metal1 880 -3060 1340 -2000 3 Cp2
port 2 e
<< end >>
