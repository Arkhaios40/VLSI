magic
tech sky130A
magscale 1 2
timestamp 1669236281
<< pwell >>
rect -1252 -10598 1252 10598
<< psubdiff >>
rect -1216 10528 1216 10562
rect -1216 10466 -1182 10528
rect 1182 10466 1216 10528
rect -1216 -10528 -1182 -10466
rect 1182 -10528 1216 -10466
rect -1216 -10562 1216 -10528
<< psubdiffcont >>
rect -1216 -10466 -1182 10466
rect 1182 -10466 1216 10466
<< xpolycontact >>
rect -1086 10000 -804 10432
rect -1086 -10432 -804 -10000
rect -708 10000 -426 10432
rect -708 -10432 -426 -10000
rect -330 10000 -48 10432
rect -330 -10432 -48 -10000
rect 48 10000 330 10432
rect 48 -10432 330 -10000
rect 426 10000 708 10432
rect 426 -10432 708 -10000
rect 804 10000 1086 10432
rect 804 -10432 1086 -10000
<< xpolyres >>
rect -1086 -10000 -804 10000
rect -708 -10000 -426 10000
rect -330 -10000 -48 10000
rect 48 -10000 330 10000
rect 426 -10000 708 10000
rect 804 -10000 1086 10000
<< locali >>
rect -1216 10528 1216 10562
rect -1216 10466 -1182 10528
rect 1182 10466 1216 10528
rect -1216 -10528 -1182 -10466
rect 1182 -10528 1216 -10466
rect -1216 -10562 1216 -10528
<< viali >>
rect -1070 10017 -820 10414
rect -692 10017 -442 10414
rect -314 10017 -64 10414
rect 64 10017 314 10414
rect 442 10017 692 10414
rect 820 10017 1070 10414
rect -1070 -10414 -820 -10017
rect -692 -10414 -442 -10017
rect -314 -10414 -64 -10017
rect 64 -10414 314 -10017
rect 442 -10414 692 -10017
rect 820 -10414 1070 -10017
<< metal1 >>
rect -1076 10414 -814 10426
rect -1076 10017 -1070 10414
rect -820 10017 -814 10414
rect -1076 10005 -814 10017
rect -698 10414 -436 10426
rect -698 10017 -692 10414
rect -442 10017 -436 10414
rect -698 10005 -436 10017
rect -320 10414 -58 10426
rect -320 10017 -314 10414
rect -64 10017 -58 10414
rect -320 10005 -58 10017
rect 58 10414 320 10426
rect 58 10017 64 10414
rect 314 10017 320 10414
rect 58 10005 320 10017
rect 436 10414 698 10426
rect 436 10017 442 10414
rect 692 10017 698 10414
rect 436 10005 698 10017
rect 814 10414 1076 10426
rect 814 10017 820 10414
rect 1070 10017 1076 10414
rect 814 10005 1076 10017
rect -1076 -10017 -814 -10005
rect -1076 -10414 -1070 -10017
rect -820 -10414 -814 -10017
rect -1076 -10426 -814 -10414
rect -698 -10017 -436 -10005
rect -698 -10414 -692 -10017
rect -442 -10414 -436 -10017
rect -698 -10426 -436 -10414
rect -320 -10017 -58 -10005
rect -320 -10414 -314 -10017
rect -64 -10414 -58 -10017
rect -320 -10426 -58 -10414
rect 58 -10017 320 -10005
rect 58 -10414 64 -10017
rect 314 -10414 320 -10017
rect 58 -10426 320 -10414
rect 436 -10017 698 -10005
rect 436 -10414 442 -10017
rect 692 -10414 698 -10017
rect 436 -10426 698 -10414
rect 814 -10017 1076 -10005
rect 814 -10414 820 -10017
rect 1070 -10414 1076 -10017
rect 814 -10426 1076 -10414
<< res1p41 >>
rect -1088 -10002 -802 10002
rect -710 -10002 -424 10002
rect -332 -10002 -46 10002
rect 46 -10002 332 10002
rect 424 -10002 710 10002
rect 802 -10002 1088 10002
<< properties >>
string FIXED_BBOX -1199 -10545 1199 10545
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 100 m 1 nx 6 wmin 1.410 lmin 0.50 rho 2000 val 142.11k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
