magic
tech sky130A
magscale 1 2
timestamp 1670987218
<< nwell >>
rect 53880 90774 56556 91408
rect 53852 84876 56528 85510
rect 53838 78808 56514 79442
rect 53924 72542 56600 73176
rect 53810 66870 56486 67504
rect 53544 60970 56220 61604
rect 53528 54972 56204 55606
rect 53346 48694 56022 49328
rect 53318 42584 55994 43218
rect 53346 36460 56022 37094
rect 53514 30786 56190 31420
rect 53628 24986 56304 25620
rect 53726 19636 56402 20270
<< metal1 >>
rect -2600 107400 2200 109200
rect 1312 104622 2846 104708
rect 1312 103188 1356 104622
rect 2790 103188 4496 104622
rect 48094 104300 48100 106100
rect 49900 104300 49906 106100
rect 1312 103116 2846 103188
rect -2600 100600 2200 102400
rect 48100 100000 49900 104300
rect 50644 103616 51073 103622
rect 53388 103616 56034 105866
rect 51073 103187 56054 103616
rect 50644 103181 51073 103187
rect 53388 103178 56054 103187
rect 55625 102572 56054 103178
rect 44494 97700 44500 99500
rect 46300 97700 46306 99500
rect 48000 98000 50000 100000
rect -2600 93800 2200 95600
rect 40694 93800 40700 95600
rect 42500 93800 42506 95600
rect 44500 94100 46300 97700
rect 53852 96518 56528 97152
rect 40700 90100 42500 93800
rect 44500 92300 49900 94100
rect 53880 90774 56556 91408
rect -2600 87000 2200 88800
rect 40700 88300 49900 90100
rect 48100 86500 49900 88300
rect 36294 83900 36300 85700
rect 38100 83900 38106 85700
rect 53852 84876 56528 85510
rect 36300 82500 38100 83900
rect -2600 80200 2200 82000
rect 36300 80700 50300 82500
rect 53838 78808 56514 79442
rect 35100 77600 36900 77606
rect 36900 75800 49700 77600
rect 35100 75794 36900 75800
rect -2600 73400 2200 75200
rect 47900 74500 49700 75800
rect 53924 72542 56600 73176
rect 35300 71000 37100 71006
rect 37100 69200 49900 71000
rect 35300 69194 37100 69200
rect -2600 66600 2200 68400
rect 48100 68100 49900 69200
rect 53810 66870 56486 67504
rect 33600 64200 35600 64400
rect 33600 62400 33700 64200
rect 35500 62400 49900 64200
rect 33600 62200 35600 62400
rect -2600 59800 2200 61600
rect 53544 60970 56220 61604
rect 33100 57400 34900 57406
rect 43500 57400 49900 58500
rect 34900 56700 49900 57400
rect 34900 55600 45300 56700
rect 33100 55594 34900 55600
rect 53528 54972 56204 55606
rect 32600 54200 34600 54400
rect -2600 52400 2200 54200
rect 32600 52400 32700 54200
rect 34500 52400 49900 54200
rect 32600 52200 34600 52400
rect 48100 50300 49900 52400
rect 53346 48694 56022 49328
rect 37600 47400 39600 47600
rect -2600 45600 2200 47400
rect 37600 45600 37700 47400
rect 39500 46100 45700 47400
rect 39500 45600 49900 46100
rect 37600 45400 39600 45600
rect 43900 44300 49900 45600
rect 53318 42584 55994 43218
rect 37800 40600 39800 40800
rect -2600 38800 2200 40600
rect 37800 38800 37900 40600
rect 39700 38800 49700 40600
rect 37800 38600 39800 38800
rect 47900 37700 49700 38800
rect 53346 36460 56022 37094
rect -2600 32000 2200 33800
rect 37200 33600 39200 33800
rect 37200 31800 37300 33600
rect 39100 31800 50100 33600
rect 37200 31600 39200 31800
rect 53514 30786 56190 31420
rect -2600 25200 2200 27000
rect 34700 26700 50500 28500
rect 34700 22800 36500 26700
rect 53628 24986 56304 25620
rect 34600 22600 36600 22800
rect 34600 20800 34700 22600
rect 36500 20800 36600 22600
rect 48300 21900 50100 23100
rect 34600 20600 36600 20800
rect -2600 18400 2200 20200
rect 37100 20100 50100 21900
rect 37100 15800 38900 20100
rect 50573 19636 50579 20270
rect 51213 19636 56402 20270
rect 37094 14000 37100 15800
rect 38900 14000 38906 15800
rect 39900 15300 50300 17100
rect -2600 11800 2200 13600
rect 39900 9200 41700 15300
rect 53880 13404 53886 13836
rect 54318 13404 57372 13836
rect 39894 7400 39900 9200
rect 41700 7400 41706 9200
rect -2600 4800 2200 6600
rect 48700 4500 50500 10900
rect 42100 2700 50500 4500
rect 42100 2400 43900 2700
rect 42094 600 42100 2400
rect 43900 600 43906 2400
<< via1 >>
rect 1356 103188 2790 104622
rect 48100 104300 49900 106100
rect 50644 103187 51073 103616
rect 44500 97700 46300 99500
rect 40700 93800 42500 95600
rect 36300 83900 38100 85700
rect 35100 75800 36900 77600
rect 35300 69200 37100 71000
rect 33700 62400 35500 64200
rect 33100 55600 34900 57400
rect 32700 52400 34500 54200
rect 37700 45600 39500 47400
rect 37900 38800 39700 40600
rect 37300 31800 39100 33600
rect 34700 20800 36500 22600
rect 50579 19636 51213 20270
rect 37100 14000 38900 15800
rect 53886 13404 54318 13836
rect 39900 7400 41700 9200
rect 42100 600 43900 2400
<< metal2 >>
rect 48100 109195 49900 109200
rect 48096 107405 48105 109195
rect 49895 107405 49904 109195
rect 48100 106100 49900 107405
rect 1270 104622 2846 104708
rect 1270 103188 1356 104622
rect 2790 103188 2846 104622
rect 48100 104294 49900 104300
rect 50649 103616 51068 103620
rect 1270 103074 2846 103188
rect 50638 103187 50644 103616
rect 51073 103187 51079 103616
rect 50649 103183 51068 103187
rect 44505 102400 46295 102404
rect 44500 102395 46300 102400
rect 44500 100605 44505 102395
rect 46295 100605 46300 102395
rect 44500 99500 46300 100605
rect 44500 97694 46300 97700
rect 40700 95600 42500 95606
rect 40700 93794 42500 93800
rect 36305 88800 38095 88804
rect 36300 88795 38100 88800
rect 36300 87005 36305 88795
rect 38095 87005 38100 88795
rect 36300 85700 38100 87005
rect 36300 83894 38100 83900
rect 35105 77600 36895 77604
rect 35094 75800 35100 77600
rect 36900 75800 36906 77600
rect 35105 75796 36895 75800
rect 35305 71000 37095 71004
rect 35294 69200 35300 71000
rect 37100 69200 37106 71000
rect 35305 69196 37095 69200
rect 33600 64200 35600 64400
rect 33600 62400 33700 64200
rect 35500 62400 35600 64200
rect 33600 62200 35600 62400
rect 33105 57400 34895 57404
rect 33094 55600 33100 57400
rect 34900 55600 34906 57400
rect 33105 55596 34895 55600
rect 32600 54200 34600 54400
rect 32600 52400 32700 54200
rect 34500 52400 34600 54200
rect 32600 52200 34600 52400
rect 37600 47400 39600 47600
rect 37600 45600 37700 47400
rect 39500 45600 39600 47400
rect 37600 45400 39600 45600
rect 37800 40600 39800 40800
rect 37800 38800 37900 40600
rect 39700 38800 39800 40600
rect 37800 38600 39800 38800
rect 37200 33600 39200 33800
rect 37200 31800 37300 33600
rect 39100 31800 39200 33600
rect 37200 31600 39200 31800
rect 34600 22600 36600 22800
rect 34600 20800 34700 22600
rect 36500 20800 36600 22600
rect 34600 20600 36600 20800
rect 50516 20270 51234 20340
rect 50516 19636 50579 20270
rect 51213 19636 51234 20270
rect 50516 19494 51234 19636
rect 37100 15800 38900 15806
rect 37100 13994 38900 14000
rect 53886 13836 54318 13842
rect 53877 13404 53886 13836
rect 54318 13404 54327 13836
rect 53886 13398 54318 13404
rect 39900 9200 41700 9206
rect 39896 7405 39900 9195
rect 41700 7405 41704 9195
rect 39900 7394 41700 7400
rect 42100 2400 43900 2406
rect 42096 605 42100 2395
rect 43900 605 43904 2395
rect 42100 594 43900 600
<< via2 >>
rect 48105 107405 49895 109195
rect 1356 103188 2790 104622
rect 50649 103192 51068 103611
rect 44505 100605 46295 102395
rect 40705 93805 42495 95595
rect 36305 87005 38095 88795
rect 35105 75805 36895 77595
rect 35305 69205 37095 70995
rect 33705 62405 35495 64195
rect 33105 55605 34895 57395
rect 32705 52405 34495 54195
rect 37705 45605 39495 47395
rect 37905 38805 39695 40595
rect 37305 31805 39095 33595
rect 34705 20805 36495 22595
rect 50579 19636 51213 20270
rect 37105 14005 38895 15795
rect 53886 13404 54318 13836
rect 39905 7405 41695 9195
rect 42105 605 43895 2395
<< metal3 >>
rect 29200 109195 49900 109200
rect 29200 107405 48105 109195
rect 49895 107405 49900 109195
rect 29200 107400 49900 107405
rect 1270 104622 2846 104708
rect -809 103188 1356 104622
rect 2790 103188 2846 104622
rect 1270 103074 2846 103188
rect 50644 103611 51073 103616
rect 50644 103192 50649 103611
rect 51068 103192 51073 103611
rect 29400 102395 46300 102400
rect 29400 100605 44505 102395
rect 46295 100605 46300 102395
rect 29400 100600 46300 100605
rect 29000 95595 42500 95600
rect 29000 93805 40705 95595
rect 42495 93805 42500 95595
rect 29000 93800 42500 93805
rect 29000 88795 38100 88800
rect 29000 87005 36305 88795
rect 38095 87005 38100 88795
rect 29000 87000 38100 87005
rect 29000 77595 36900 77600
rect 29000 75805 35105 77595
rect 36895 75805 36900 77595
rect 29000 75800 36900 75805
rect 29200 70995 37100 71000
rect 29200 69205 35305 70995
rect 37095 69205 37100 70995
rect 29200 69200 37100 69205
rect 33600 64200 35600 64400
rect 28800 64195 35600 64200
rect 28800 62405 33705 64195
rect 35495 62405 35600 64195
rect 28800 62400 35600 62405
rect 33600 62200 35600 62400
rect 28000 57395 34900 57400
rect 28000 55605 33105 57395
rect 34895 55605 34900 57395
rect 28000 55600 34900 55605
rect 32600 54200 34600 54400
rect 29400 54195 34600 54200
rect 29400 52405 32705 54195
rect 34495 52405 34600 54195
rect 29400 52400 34600 52405
rect 32600 52200 34600 52400
rect 37600 47400 39600 47600
rect 29200 47395 39600 47400
rect 29200 45605 37705 47395
rect 39495 45605 39600 47395
rect 29200 45600 39600 45605
rect 37600 45400 39600 45600
rect 37800 40600 39800 40800
rect 29000 40595 39800 40600
rect 29000 38805 37905 40595
rect 39695 38805 39800 40595
rect 29000 38800 39800 38805
rect 37800 38600 39800 38800
rect 37200 33600 39200 33800
rect 29000 33595 39200 33600
rect 29000 31805 37305 33595
rect 39095 31805 39200 33595
rect 29000 31800 39200 31805
rect 37200 31600 39200 31800
rect 34600 22600 36600 22800
rect 29000 22595 36600 22600
rect 29000 20805 34705 22595
rect 36495 20805 36600 22595
rect 29000 20800 36600 20805
rect 34600 20600 36600 20800
rect 50644 20275 51073 103192
rect 50574 20270 51218 20275
rect 50574 19636 50579 20270
rect 51213 19636 51218 20270
rect 50574 19631 51218 19636
rect 29000 15795 38900 15800
rect 29000 14005 37105 15795
rect 38895 14005 38900 15795
rect 29000 14000 38900 14005
rect 50644 13836 51073 19631
rect 53881 13836 54323 13841
rect 50478 13404 53886 13836
rect 54318 13404 54323 13836
rect 53881 13399 54323 13404
rect 28800 9195 41700 9200
rect 28800 7405 39905 9195
rect 41695 7405 41700 9195
rect 28800 7400 41700 7405
rect 27800 2395 43900 2400
rect 27800 605 42105 2395
rect 43895 605 43900 2395
rect 27800 600 43900 605
<< metal4 >>
rect 93200 97800 106200 100200
rect 93200 91600 106200 94000
rect 93200 86000 106200 88400
rect 93200 80200 106200 82600
rect 93200 74200 106200 76600
rect 93200 67400 106200 69800
rect 93200 62000 106200 64400
rect 93200 57400 106200 59800
rect 67000 50400 106200 52800
rect 79200 44200 106200 46400
rect 80200 38000 106200 40400
rect 81000 32000 106200 34400
rect 81600 26000 106200 28600
rect 83400 20000 106200 22600
rect 85000 14800 106200 17400
rect 87000 8400 106200 11000
use NMOSR2Stg1  NMOSR2Stg1_0
timestamp 1670983913
transform 1 0 3040 0 1 55508
box -3040 -508 28369 53400
use NMOSR2Stg1  NMOSR2Stg1_1
timestamp 1670983913
transform 1 0 3040 0 1 508
box -3040 -508 28369 53400
use PMOSOutStg  PMOSOutStg_0
timestamp 1670438645
transform 1 0 54188 0 1 15326
box -6188 -8326 49583 89584
<< labels >>
rlabel metal1 -2600 107400 2200 109200 7 IN_X0_I+
port 0 w
rlabel metal4 93200 97800 106200 100200 3 OUT_Y0_I+
port 1 e
rlabel metal1 -2600 100600 2200 102400 7 IN_X0_I-
port 2 w
rlabel metal4 93200 91600 106200 94000 3 OUT_Y0_I-
port 3 e
rlabel metal1 -2600 93800 2200 95600 7 IN_X0_Q+
port 4 w
rlabel metal4 93200 86000 106200 88400 3 OUT_X0_Q+
port 5 e
rlabel metal1 -2600 87000 2200 88800 7 IN_X0_Q-
port 6 w
rlabel metal4 93200 80200 106200 82600 3 OUT_X0_Q-
port 7 e
rlabel metal1 -2600 80200 2200 82000 7 IN_X2_I+
port 8 w
rlabel metal4 93200 74200 106200 76600 3 OUT_Y1_I+
port 9 e
rlabel metal1 -2600 73400 2200 75200 7 IN_X2_I-
port 10 w
rlabel metal1 -2600 66600 2200 68400 7 IN_X2_Q+
port 12 w
rlabel metal4 93200 62000 106200 64400 3 OUT_Y1_Q+
port 13 e
rlabel metal4 93200 67400 106200 69800 3 OUT_Y1_I-
port 11 e
rlabel metal1 -2600 59800 2200 61600 7 IN_X2_Q-
port 14 w
rlabel metal4 93200 57400 106200 59800 3 OUT_Y1_Q-
port 15 e
rlabel metal1 -2600 52400 2200 54200 7 IN_X1_I+
port 16 w
rlabel metal1 -2600 45600 2200 47400 7 IN_X1_I-
port 18 w
rlabel metal1 -2600 38800 2200 40600 7 IN_X1_Q+
port 20 w
rlabel metal1 -2600 32000 2200 33800 7 IN_X1_Q-
port 22 w
rlabel metal1 -2600 25200 2200 27000 7 IN_X3_I+
port 24 w
rlabel metal1 -2600 18400 2200 20200 7 IN_X3_I-
port 26 w
rlabel metal1 -2600 11800 2200 13600 7 IN_X3_Q+
port 28 w
rlabel metal1 -2600 4800 2200 6600 7 IN_X3_Q-
port 30 w
rlabel metal4 67000 50400 106200 52800 3 OUT_Y2_I+
port 17 e
rlabel metal4 79200 44200 106200 46400 3 OUT_Y2_I-
port 19 e
rlabel metal4 80200 38000 106200 40400 3 OUT_Y2_Q+
port 21 e
rlabel metal4 81000 32000 106200 34400 3 OUT_Y2_Q-
port 23 e
rlabel metal4 81600 26000 106200 28600 3 OUT_Y3_I+
port 25 e
rlabel metal4 83400 20000 106200 22600 3 OUT_Y3_I-
port 27 e
rlabel metal4 85000 14800 106200 17400 3 OUT_Y3_Q+
port 29 e
rlabel metal4 87000 8400 106200 11000 3 OUT_Y3_Q-
port 31 e
rlabel metal1 53388 103178 56034 105866 1 VDD!
port 32 n
<< end >>
