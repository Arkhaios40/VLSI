magic
tech sky130A
magscale 1 2
timestamp 1669545529
<< pwell >>
rect -400 8400 456 16854
<< mvnmos >>
rect -172 8658 228 16658
<< mvndiff >>
rect -230 16646 -172 16658
rect -230 8670 -218 16646
rect -184 8670 -172 16646
rect -230 8658 -172 8670
rect 228 16646 286 16658
rect 228 8670 240 16646
rect 274 8670 286 16646
rect 228 8658 286 8670
<< mvndiffc >>
rect -218 8670 -184 16646
rect 240 8670 274 16646
<< mvpsubdiff >>
rect -364 16760 420 16818
rect -364 16710 -306 16760
rect -364 8544 -352 16710
rect -318 8544 -306 16710
rect 362 16710 420 16760
rect -364 8494 -306 8544
rect 362 8544 374 16710
rect 408 8544 420 16710
rect 362 8494 420 8544
rect -364 8436 420 8494
<< mvpsubdiffcont >>
rect -352 8544 -318 16710
rect 374 8544 408 16710
<< poly >>
rect -172 16658 228 16684
rect -172 8620 228 8658
rect -172 8586 -156 8620
rect 212 8586 228 8620
rect -172 8570 228 8586
<< polycont >>
rect -156 8586 212 8620
<< locali >>
rect -352 16772 408 16806
rect -352 16710 -318 16772
rect 374 16710 408 16772
rect -218 16646 -184 16662
rect -218 8654 -184 8670
rect 240 16646 274 16662
rect 240 8654 274 8670
rect -172 8586 -156 8620
rect 212 8586 228 8620
rect -352 8520 -318 8544
rect 374 8520 408 8544
<< viali >>
rect -218 8670 -184 16646
rect 240 8670 274 16646
rect -156 8586 212 8620
<< metal1 >>
rect -224 16646 -178 16658
rect -224 8670 -218 16646
rect -184 8670 -178 16646
rect -224 8658 -178 8670
rect 234 16646 280 16658
rect 234 8670 240 16646
rect 274 8670 280 16646
rect 234 8658 280 8670
rect -168 8620 224 8626
rect -168 8586 -156 8620
rect 212 8586 224 8620
rect -168 8580 224 8586
<< metal2 >>
rect -1340 8680 -940 16640
rect 1860 8680 2262 16640
rect -1329 7951 -589 8290
rect 1548 7952 2288 8289
rect -1340 7400 -240 7760
rect 1549 7015 2285 7305
use sky130_fd_pr__nfet_g5v0d10v5_UBJTTH  sky130_fd_pr__nfet_g5v0d10v5_UBJTTH_0
timestamp 1669545529
transform -1 0 888 0 -1 12627
box -1400 -4227 2228 5633
<< labels >>
rlabel metal2 -1340 8680 -940 16640 7 D_Pin_L
port 0 w
rlabel metal2 1860 8680 2262 16640 3 D_Pin_R
port 1 e
rlabel metal2 -1329 7951 -589 8290 7 D_In_L
port 2 w
rlabel metal2 1548 7952 2288 8289 3 D_In_R
port 3 e
rlabel metal2 -1340 7400 -240 7760 7 NMOS_Vs
port 4 w
rlabel metal2 1549 7015 2285 7305 3 Body
port 5 e
<< end >>
