** sch_path: /home/arkhaios/Project/xschem/PrimalStructures/CurRefResistor.sch
**.subckt CurRefResistor Pin1 Pin2
*.iopin Pin1
*.iopin Pin2
XR1 Pin2 Pin1 GND sky130_fd_pr__res_xhigh_po_1p41 L=40 mult=1 m=1
**.ends
.GLOBAL GND
.end
