magic
tech sky130A
magscale 1 2
timestamp 1669614457
<< locali >>
rect -77 18137 455 18156
rect -77 17692 -47 18137
rect 429 17692 455 18137
rect -77 17072 455 17692
rect 7912 17178 8637 17652
rect -8596 16770 -5270 16776
rect -8596 16118 -8590 16770
rect -7938 16118 -5270 16770
rect -8596 16112 -5270 16118
rect 1526 16662 2940 16668
rect 1526 16006 1532 16662
rect 2188 16006 2940 16662
rect 1526 16000 2940 16006
<< viali >>
rect -47 17692 429 18137
rect 7912 17652 8637 18377
rect -8590 16118 -7938 16770
rect 1532 16006 2188 16662
<< metal1 >>
rect -32934 19943 -30724 19960
rect -23393 19943 -22680 19960
rect -16468 19943 19446 19960
rect -34107 18377 19446 19943
rect -34107 18137 7912 18377
rect -34107 17692 -47 18137
rect 429 17692 7912 18137
rect -34107 17652 7912 17692
rect 8637 17652 19446 18377
rect -34107 17645 19446 17652
rect -34107 -2661 -33393 17645
rect -32934 17644 -30724 17645
rect -30058 15498 -29232 17645
rect -21522 15492 -20690 17645
rect -16468 17644 19446 17645
rect -3247 16968 -2809 17644
rect 3769 17050 4207 17644
rect -9914 16776 -9250 16782
rect -9250 16770 -7926 16776
rect -9250 16118 -8590 16770
rect -7938 16118 -7926 16770
rect -9250 16112 -7926 16118
rect 1526 16662 2194 16674
rect -9914 16106 -9250 16112
rect 1526 16006 1532 16662
rect 2188 16006 2194 16662
rect 13478 16629 14533 17644
rect 1526 15994 2194 16006
rect 1528 15684 2192 15994
rect 1522 15020 1528 15684
rect 2192 15020 2198 15684
rect 13472 15574 13478 16629
rect 14533 15574 14539 16629
rect -6994 13942 -6594 13948
rect -6594 13542 -5544 13942
rect 1509 13683 1515 14085
rect 1917 13683 2571 14085
rect -6994 13536 -6594 13542
rect -29774 8032 -29110 8956
rect -19823 7635 -19165 9149
rect -4314 8948 -3594 11088
rect 3948 8948 4668 8954
rect -4314 8228 3948 8948
rect 3948 8222 4668 8228
rect 5399 8895 6129 11209
rect 7168 8895 7898 8901
rect 5399 8165 7168 8895
rect 7168 8159 7898 8165
rect -29774 7362 -29110 7368
rect -19829 6977 -19823 7635
rect -19165 6977 -19159 7635
rect -34109 -3379 -31763 -2661
rect -9917 -12560 -9327 -9878
rect -930 -11574 -924 -11290
rect -640 -11574 -634 -11290
rect -924 -12560 -640 -11574
rect 6502 -11675 6508 -11177
rect 7006 -11675 7012 -11177
rect 6508 -12560 7006 -11675
rect -33596 -13005 18784 -12560
rect -33596 -13595 -22188 -13005
rect -21598 -13595 18784 -13005
rect -33596 -14876 18784 -13595
<< via1 >>
rect -9914 16112 -9250 16776
rect 1528 15020 2192 15684
rect 13478 15574 14533 16629
rect -6994 13542 -6594 13942
rect 1515 13683 1917 14085
rect -29774 7368 -29110 8032
rect 3948 8228 4668 8948
rect 7168 8165 7898 8895
rect -19823 6977 -19165 7635
rect -924 -11574 -640 -11290
rect 6508 -11675 7006 -11177
rect -22188 -13595 -21598 -13005
<< metal2 >>
rect -9920 16112 -9914 16776
rect -9250 16112 -9244 16776
rect 13478 16629 14533 16635
rect -9914 15679 -9250 16112
rect 221 15684 875 15688
rect 1528 15684 2192 15690
rect -9914 15025 -9909 15679
rect -9255 15025 -9250 15679
rect -9914 15020 -9250 15025
rect 216 15679 1528 15684
rect 216 15025 221 15679
rect 875 15025 1528 15679
rect 216 15020 1528 15025
rect -9909 15016 -9255 15020
rect 221 15016 875 15020
rect 1528 15014 2192 15020
rect 1515 14085 1917 14091
rect -11668 13542 -6994 13942
rect -6594 13542 -6588 13942
rect -11668 9314 -11268 13542
rect 1515 10141 1917 13683
rect -8468 9739 1917 10141
rect -8468 9313 -8066 9739
rect 3942 8228 3948 8948
rect 4668 8228 4674 8948
rect -29780 7368 -29774 8032
rect -28520 7368 -28511 8032
rect -19823 7635 -19165 7641
rect -19823 1531 -19165 6977
rect 3948 3704 4668 8228
rect 7162 8165 7168 8895
rect 7898 8165 7904 8895
rect 7168 3674 7898 8165
rect 8675 8067 9334 8072
rect 8671 7418 8680 8067
rect 9329 7418 9338 8067
rect 13478 7644 14533 15574
rect 8675 2709 9334 7418
rect -19823 873 -16767 1531
rect -11649 1141 -11640 1480
rect -11301 1141 -11292 1480
rect -8420 1142 -8411 1479
rect -8074 1142 -8065 1479
rect -17425 -1384 -16767 873
rect -17425 -2040 -12354 -1384
rect -17425 -2041 -16767 -2040
rect -13010 -2930 -12354 -2040
rect -11592 -2608 -11232 950
rect -8333 -1373 -8043 495
rect 18925 389 18934 709
rect 19254 389 19263 709
rect -8333 -1663 -637 -1373
rect -11592 -2968 -6552 -2608
rect -924 -11290 -640 -1663
rect -924 -11580 -640 -11574
rect 6508 -11177 7006 -4862
rect -22188 -13005 -21598 -11650
rect 6508 -11681 7006 -11675
rect -22194 -13595 -22188 -13005
rect -21598 -13595 -21592 -13005
<< via2 >>
rect -9909 15025 -9255 15679
rect 221 15025 875 15679
rect -29184 7368 -29110 8032
rect -29110 7368 -28520 8032
rect 8680 7418 9329 8067
rect -11640 1141 -11301 1480
rect -8411 1142 -8074 1479
rect 18934 389 19254 709
<< metal3 >>
rect -14622 15679 9336 15684
rect -14622 15025 -9909 15679
rect -9255 15025 221 15679
rect 875 15025 9336 15679
rect -14622 15020 9336 15025
rect -14622 13414 -13958 15020
rect -17118 12750 -13958 13414
rect -17118 8062 -16454 12750
rect -29189 8032 -28515 8037
rect -27077 8032 -16454 8062
rect -29189 7368 -29184 8032
rect -28520 7403 -16454 8032
rect 8675 8067 9334 15020
rect 8675 7418 8680 8067
rect 9329 7418 9334 8067
rect 8675 7413 9334 7418
rect -28520 7368 -26595 7403
rect -29189 7363 -28515 7368
rect -24108 -886 -23444 7403
rect -11645 1480 -11296 1485
rect -12723 1141 -12717 1480
rect -12378 1141 -11640 1480
rect -11301 1141 -11296 1480
rect -11645 1136 -11296 1141
rect -8416 1479 -8069 1484
rect -8416 1142 -8411 1479
rect -8074 1142 -7493 1479
rect -7156 1142 -7150 1479
rect -8416 1137 -8069 1142
rect 18929 709 19259 714
rect 18929 389 18934 709
rect 19254 389 20560 709
rect 20880 389 20886 709
rect 18929 384 19259 389
rect -19166 -886 -18374 -870
rect -24108 -1550 -18374 -886
rect -19166 -1636 -18374 -1550
<< via3 >>
rect -12717 1141 -12378 1480
rect -7493 1142 -7156 1479
rect 20560 389 20880 709
<< metal4 >>
rect -12718 1480 -12377 1481
rect -13368 1141 -12717 1480
rect -12378 1141 -12377 1480
rect -7494 1479 -7155 1480
rect -7494 1142 -7493 1479
rect -7156 1142 -6357 1479
rect -7494 1141 -7155 1142
rect -12718 1140 -12377 1141
rect 20559 709 20881 710
rect 20559 389 20560 709
rect 20880 389 22594 709
rect 20559 388 20881 389
<< via4 >>
rect -13707 1141 -13368 1480
rect -6357 1142 -6020 1479
rect 22594 389 22914 709
<< metal5 >>
rect -13731 1480 -13344 1504
rect -14899 1479 -13707 1480
rect -37866 1142 -13707 1479
rect -14899 1141 -13707 1142
rect -13368 1141 -13344 1480
rect -13731 1117 -13344 1141
rect -6381 1479 -5996 1503
rect -6381 1142 -6357 1479
rect -6020 1142 -5996 1479
rect -6381 1118 -5996 1142
rect -6356 169 -6019 1118
rect 22570 709 22938 733
rect 22570 389 22594 709
rect 22914 389 27270 709
rect 22570 365 22938 389
rect -37954 -168 -6019 169
use ConnectedNMOSPair  ConnectedNMOSPair_0
timestamp 1669244576
transform 1 0 -7172 0 1 -10384
box -5846 -84 5646 8110
use ConnectedPMOSPair  ConnectedPMOSPair_1
timestamp 1669614457
transform 1 0 -22909 0 1 9557
box -8826 -1262 8104 7824
use CurrentRef  CurrentRef_0
timestamp 1669422754
transform 1 0 -24709 0 1 -14875
box -7985 2635 11290 22119
use DifferentialPair  DifferentialPair_0
timestamp 1669545529
transform 1 0 -10328 0 1 -6810
box -1340 6994 2288 16854
use GainStage  GainStage_0
timestamp 1669543272
transform 1 0 7158 0 1 509
box -4840 -5869 12280 8287
use PMOSPair  PMOSPair_0
timestamp 1669589303
transform 1 0 -5026 0 1 9364
box -848 1666 6432 8042
use PMOSPair  PMOSPair_1
timestamp 1669589303
transform 1 0 3166 0 1 9446
box -848 1666 6432 8042
<< labels >>
rlabel metal1 -34107 17645 -4742 19943 1 VDD
port 0 n
rlabel metal5 -37866 1142 -13707 1479 7 In+
port 1 w
rlabel metal5 -37954 -168 -6019 169 7 In-
port 2 w
rlabel space 0 0 0 0 3 Out
rlabel metal5 22914 389 27270 709 3 Out
port 3 e
rlabel metal1 -33596 -14876 -22188 -12560 5 Ground
port 4 s
<< end >>
