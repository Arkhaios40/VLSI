magic
tech sky130A
magscale 1 2
timestamp 1669425766
<< pwell >>
rect -428 -4305 428 4305
<< mvnmos >>
rect -200 47 200 4047
rect -200 -4109 200 -109
<< mvndiff >>
rect -258 4035 -200 4047
rect -258 59 -246 4035
rect -212 59 -200 4035
rect -258 47 -200 59
rect 200 4035 258 4047
rect 200 59 212 4035
rect 246 59 258 4035
rect 200 47 258 59
rect -258 -121 -200 -109
rect -258 -4097 -246 -121
rect -212 -4097 -200 -121
rect -258 -4109 -200 -4097
rect 200 -121 258 -109
rect 200 -4097 212 -121
rect 246 -4097 258 -121
rect 200 -4109 258 -4097
<< mvndiffc >>
rect -246 59 -212 4035
rect 212 59 246 4035
rect -246 -4097 -212 -121
rect 212 -4097 246 -121
<< mvpsubdiff >>
rect -392 4211 392 4269
rect -392 4161 -334 4211
rect -392 -4161 -380 4161
rect -346 -4161 -334 4161
rect 334 4161 392 4211
rect -392 -4211 -334 -4161
rect 334 -4161 346 4161
rect 380 -4161 392 4161
rect 334 -4211 392 -4161
rect -392 -4269 392 -4211
<< mvpsubdiffcont >>
rect -380 -4161 -346 4161
rect 346 -4161 380 4161
<< poly >>
rect -200 4119 200 4135
rect -200 4085 -184 4119
rect 184 4085 200 4119
rect -200 4047 200 4085
rect -200 21 200 47
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect -200 -4135 200 -4109
<< polycont >>
rect -184 4085 184 4119
rect -184 -71 184 -37
<< locali >>
rect -380 4223 380 4257
rect -380 4161 -346 4223
rect 346 4161 380 4223
rect -200 4085 -184 4119
rect 184 4085 200 4119
rect -246 4035 -212 4051
rect -246 43 -212 59
rect 212 4035 246 4051
rect 212 43 246 59
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -121 -212 -105
rect -246 -4113 -212 -4097
rect 212 -121 246 -105
rect 212 -4113 246 -4097
rect -380 -4223 -346 -4161
rect 346 -4223 380 -4161
rect -380 -4257 380 -4223
<< viali >>
rect -184 4085 184 4119
rect -246 59 -212 4035
rect 212 59 246 4035
rect -184 -71 184 -37
rect -246 -4097 -212 -121
rect 212 -4097 246 -121
<< metal1 >>
rect -196 4119 196 4125
rect -196 4085 -184 4119
rect 184 4085 196 4119
rect -196 4079 196 4085
rect -252 4035 -206 4047
rect -252 59 -246 4035
rect -212 59 -206 4035
rect -252 47 -206 59
rect 206 4035 252 4047
rect 206 59 212 4035
rect 246 59 252 4035
rect 206 47 252 59
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -121 -206 -109
rect -252 -4097 -246 -121
rect -212 -4097 -206 -121
rect -252 -4109 -206 -4097
rect 206 -121 252 -109
rect 206 -4097 212 -121
rect 246 -4097 252 -121
rect 206 -4109 252 -4097
<< properties >>
string FIXED_BBOX -363 -4240 363 4240
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 20 l 2 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
