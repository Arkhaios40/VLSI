magic
tech sky130A
magscale 1 2
timestamp 1669589303
<< locali >>
rect -398 7576 -212 7578
rect -398 6612 84 7576
rect -398 6086 -212 6612
rect 8 6252 4646 6454
rect -398 5718 92 6086
rect -398 5188 -212 5718
rect 4476 5562 4646 6252
rect 0 5348 4646 5562
rect -398 4820 80 5188
rect -398 4280 -212 4820
rect 4476 4660 4646 5348
rect 0 4446 4646 4660
rect -398 3912 70 4280
rect -398 3370 -212 3912
rect 4476 3752 4646 4446
rect -4 3538 4646 3752
rect -398 3002 70 3370
rect -398 2486 -212 3002
rect 4476 2850 4646 3538
rect -18 2636 4646 2850
rect 4476 2574 4646 2636
rect -398 2104 74 2486
<< metal1 >>
rect 198 7604 6084 8042
rect -848 6466 -476 6576
rect 184 6466 4062 6580
rect -848 6206 4062 6466
rect -848 4680 -476 6206
rect 184 6102 4062 6206
rect 180 5560 4058 5694
rect 4676 5560 4984 5634
rect 180 5344 4984 5560
rect 180 5216 4058 5344
rect 168 4680 4006 4780
rect -848 4420 4006 4680
rect -848 2878 -476 4420
rect 168 4318 4006 4420
rect 162 3746 4040 3876
rect 4676 3746 4984 5344
rect 162 3530 4984 3746
rect 162 3398 4040 3530
rect 188 2878 4026 2978
rect -848 2618 4026 2878
rect -848 2542 -476 2618
rect 188 2516 4026 2618
rect 182 1932 4048 2086
rect 4676 1932 4984 3530
rect 182 1670 4984 1932
rect 182 1668 4916 1670
rect 4398 1666 4916 1668
use sky130_fd_pr__pfet_g5v0d10v5_97TZA6  XM7
timestamp 1668107812
transform 0 -1 2139 1 0 5900
box -458 -2297 458 2297
use sky130_fd_pr__pfet_g5v0d10v5_97TZA6  XM8
timestamp 1668107812
transform 0 -1 2133 1 0 5004
box -458 -2297 458 2297
use sky130_fd_pr__pfet_g5v0d10v5_97TZA6  XM9
timestamp 1668107812
transform 0 -1 2121 1 0 4092
box -458 -2297 458 2297
use sky130_fd_pr__pfet_g5v0d10v5_97TZA6  XM10
timestamp 1668107812
transform 0 -1 2117 1 0 3188
box -458 -2297 458 2297
use sky130_fd_pr__pfet_g5v0d10v5_97TZA6  XM11
timestamp 1668107812
transform 0 -1 2113 1 0 2296
box -458 -2297 458 2297
use sky130_fd_pr__pfet_g5v0d10v5_97BMAW  XM12
timestamp 1668639803
transform 0 1 3135 -1 0 7100
box -758 -3297 758 3297
<< labels >>
rlabel metal1 322 7900 3470 8008 1 Vs
port 0 n
rlabel locali 4506 5724 4626 6228 3 body
port 1 e
rlabel metal1 -804 5544 -638 6472 7 CenterTap
port 2 w
rlabel locali -356 6812 -254 7362 7 Vp
port 3 w
rlabel space 182 1668 4048 2090 5 Vd
port 5 s
<< end >>
