magic
tech sky130A
magscale 1 2
timestamp 1669244576
<< locali >>
rect -2762 6244 -2434 6260
rect -2762 5910 -2218 6244
rect -2762 5398 -2434 5910
rect 2134 5724 2342 6470
rect -2270 5580 2342 5724
rect -2762 5064 -2208 5398
rect -2762 4538 -2434 5064
rect 2134 4868 2342 5580
rect -2270 4724 2342 4868
rect -2762 4204 -2218 4538
rect -2762 3680 -2434 4204
rect 2134 4016 2342 4724
rect -2284 3872 2342 4016
rect -2762 3346 -2220 3680
rect -2762 2826 -2434 3346
rect 2134 3160 2342 3872
rect -2278 3016 2342 3160
rect -2762 2492 -2218 2826
rect -2762 1968 -2434 2492
rect 2134 2330 2342 3016
rect -2312 2130 2342 2330
rect -2312 2128 2326 2130
rect -2762 1872 -2206 1968
rect -2758 1030 -2206 1872
<< metal1 >>
rect -3026 5780 -2370 6752
rect 2376 6750 2612 6762
rect 852 6540 2612 6750
rect -2128 6486 2612 6540
rect -2128 6276 1740 6486
rect -2082 5780 1726 5878
rect -3034 5516 1726 5780
rect -3026 4088 -2370 5516
rect -2082 5426 1726 5516
rect -2114 4928 1680 5008
rect 2376 4928 2612 6486
rect -2114 4680 2612 4928
rect -2114 4570 1680 4680
rect -2100 4088 1708 4166
rect -3026 3824 1708 4088
rect -3026 2384 -2370 3824
rect -2100 3714 1708 3824
rect -2132 3218 1662 3310
rect 2376 3218 2612 4680
rect -2132 2970 2612 3218
rect -2132 2872 1662 2970
rect 2376 2954 2612 2970
rect -2114 2430 -326 2448
rect -2178 2384 -326 2430
rect -3026 2088 -326 2384
rect -3026 1998 -2370 2088
rect -2114 2004 -326 2088
rect -2100 22 -234 1016
use sky130_fd_pr__nfet_g5v0d10v5_HYQESV  sky130_fd_pr__nfet_g5v0d10v5_HYQESV_0
timestamp 1668098548
transform 0 -1 -209 1 0 6077
box -428 -2227 428 2227
use sky130_fd_pr__nfet_g5v0d10v5_HYQESV  sky130_fd_pr__nfet_g5v0d10v5_HYQESV_1
timestamp 1668098548
transform 0 -1 -209 1 0 2662
box -428 -2227 428 2227
use sky130_fd_pr__nfet_g5v0d10v5_HYQESV  sky130_fd_pr__nfet_g5v0d10v5_HYQESV_2
timestamp 1668098548
transform 0 -1 -211 1 0 3513
box -428 -2227 428 2227
use sky130_fd_pr__nfet_g5v0d10v5_HYQESV  sky130_fd_pr__nfet_g5v0d10v5_HYQESV_3
timestamp 1668098548
transform 0 -1 -212 1 0 4369
box -428 -2227 428 2227
use sky130_fd_pr__nfet_g5v0d10v5_HYQESV  sky130_fd_pr__nfet_g5v0d10v5_HYQESV_4
timestamp 1668098548
transform 0 -1 -209 1 0 5223
box -428 -2227 428 2227
use sky130_fd_pr__nfet_g5v0d10v5_VSVLYK  sky130_fd_pr__nfet_g5v0d10v5_VSVLYK_0
timestamp 1668623350
transform 0 -1 -1203 1 0 1500
box -728 -1227 728 1227
<< labels >>
rlabel metal1 -2855 2839 -2396 6731 1 exists
rlabel metal1 -406 670 -308 762 5 S
port 3 s
rlabel locali 2162 6180 2258 6308 1 Vnbody
port 2 n
rlabel locali -2686 1674 -2600 1782 7 Vn
port 1 w
rlabel metal1 -2734 6520 -2638 6648 1 Vd
port 0 n
<< end >>
