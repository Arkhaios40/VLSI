magic
tech sky130A
magscale 1 2
timestamp 1670361013
<< nwell >>
rect -1458 -597 1458 597
<< mvpmos >>
rect -1200 -300 1200 300
<< mvpdiff >>
rect -1258 288 -1200 300
rect -1258 -288 -1246 288
rect -1212 -288 -1200 288
rect -1258 -300 -1200 -288
rect 1200 288 1258 300
rect 1200 -288 1212 288
rect 1246 -288 1258 288
rect 1200 -300 1258 -288
<< mvpdiffc >>
rect -1246 -288 -1212 288
rect 1212 -288 1246 288
<< mvnsubdiff >>
rect -1392 519 1392 531
rect -1392 485 -1284 519
rect 1284 485 1392 519
rect -1392 473 1392 485
rect -1392 423 -1334 473
rect -1392 -423 -1380 423
rect -1346 -423 -1334 423
rect 1334 423 1392 473
rect -1392 -473 -1334 -423
rect 1334 -423 1346 423
rect 1380 -423 1392 423
rect 1334 -473 1392 -423
rect -1392 -485 1392 -473
rect -1392 -519 -1284 -485
rect 1284 -519 1392 -485
rect -1392 -531 1392 -519
<< mvnsubdiffcont >>
rect -1284 485 1284 519
rect -1380 -423 -1346 423
rect 1346 -423 1380 423
rect -1284 -519 1284 -485
<< poly >>
rect -1200 381 1200 397
rect -1200 347 -1184 381
rect 1184 347 1200 381
rect -1200 300 1200 347
rect -1200 -347 1200 -300
rect -1200 -381 -1184 -347
rect 1184 -381 1200 -347
rect -1200 -397 1200 -381
<< polycont >>
rect -1184 347 1184 381
rect -1184 -381 1184 -347
<< locali >>
rect -1380 485 -1284 519
rect 1284 485 1380 519
rect -1380 423 -1346 485
rect 1346 423 1380 485
rect -1200 347 -1184 381
rect 1184 347 1200 381
rect -1246 288 -1212 304
rect -1246 -304 -1212 -288
rect 1212 288 1246 304
rect 1212 -304 1246 -288
rect -1200 -381 -1184 -347
rect 1184 -381 1200 -347
rect -1380 -485 -1346 -423
rect 1346 -485 1380 -423
rect -1380 -519 -1284 -485
rect 1284 -519 1380 -485
<< viali >>
rect -1184 347 1184 381
rect -1246 -288 -1212 288
rect 1212 -288 1246 288
rect -1184 -381 1184 -347
<< metal1 >>
rect -1196 381 1196 387
rect -1196 347 -1184 381
rect 1184 347 1196 381
rect -1196 341 1196 347
rect -1252 288 -1206 300
rect -1252 -288 -1246 288
rect -1212 -288 -1206 288
rect -1252 -300 -1206 -288
rect 1206 288 1252 300
rect 1206 -288 1212 288
rect 1246 -288 1252 288
rect 1206 -300 1252 -288
rect -1196 -347 1196 -341
rect -1196 -381 -1184 -347
rect 1184 -381 1196 -347
rect -1196 -387 1196 -381
<< properties >>
string FIXED_BBOX -1363 -502 1363 502
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 3 l 12 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
