magic
tech sky130A
magscale 1 2
timestamp 1669545529
<< pwell >>
rect -428 -4227 428 4227
<< mvnmos >>
rect -200 -4031 200 3969
<< mvndiff >>
rect -258 3957 -200 3969
rect -258 -4019 -246 3957
rect -212 -4019 -200 3957
rect -258 -4031 -200 -4019
rect 200 3957 258 3969
rect 200 -4019 212 3957
rect 246 -4019 258 3957
rect 200 -4031 258 -4019
<< mvndiffc >>
rect -246 -4019 -212 3957
rect 212 -4019 246 3957
<< mvpsubdiff >>
rect -392 4133 392 4191
rect -392 4083 -334 4133
rect -392 -4083 -380 4083
rect -346 -4083 -334 4083
rect 334 4083 392 4133
rect -392 -4133 -334 -4083
rect 334 -4083 346 4083
rect 380 -4083 392 4083
rect 334 -4133 392 -4083
rect -392 -4191 392 -4133
<< mvpsubdiffcont >>
rect -380 -4083 -346 4083
rect 346 -4083 380 4083
<< poly >>
rect -200 4041 200 4057
rect -200 4007 -184 4041
rect 184 4007 200 4041
rect -200 3969 200 4007
rect -200 -4057 200 -4031
<< polycont >>
rect -184 4007 184 4041
<< locali >>
rect 228 5307 528 5627
rect 167 4337 168 4407
rect -380 4083 -346 4107
rect -172 4041 168 4337
rect 328 4083 528 5307
rect -200 4007 -184 4041
rect 184 4007 200 4041
rect -246 3957 -212 3973
rect -246 -4035 -212 -4019
rect 212 3957 246 3973
rect 212 -4035 246 -4019
rect 328 -4033 346 4083
rect -380 -4145 -346 -4083
rect 380 -4033 528 4083
rect 688 4007 1028 4337
rect 346 -4145 380 -4083
rect -380 -4179 380 -4145
<< viali >>
rect -92 5307 228 5627
rect -172 4337 167 4676
rect -184 4007 184 4041
rect -246 -4019 -212 3957
rect 212 -4019 246 3957
rect 688 4337 1028 4677
<< metal1 >>
rect -104 5627 240 5633
rect -104 5616 -92 5627
rect -667 5317 -661 5616
rect -362 5317 -92 5616
rect -104 5307 -92 5317
rect 228 5307 240 5627
rect -104 5301 240 5307
rect 288 4867 768 5227
rect 1128 4867 1134 5227
rect -184 4676 179 4682
rect -184 4675 -172 4676
rect -666 4338 -660 4675
rect -323 4338 -172 4675
rect -184 4337 -172 4338
rect 167 4337 179 4676
rect -184 4331 179 4337
rect -196 4041 196 4047
rect -196 4007 -184 4041
rect 184 4007 196 4041
rect -196 4001 196 4007
rect -252 3957 -206 3969
rect -252 3947 -246 3957
rect -1012 3907 -246 3947
rect -1012 -3973 -972 3907
rect -612 -3973 -246 3907
rect -1012 -4013 -246 -3973
rect -252 -4019 -246 -4013
rect -212 -4019 -206 3957
rect -252 -4031 -206 -4019
rect 206 3957 252 3969
rect 206 -4019 212 3957
rect 246 3947 252 3957
rect 288 3947 568 4867
rect 682 4677 1034 4689
rect 682 4337 688 4677
rect 1028 4676 1034 4677
rect 1028 4337 1138 4676
rect 1477 4337 1483 4676
rect 682 4325 1034 4337
rect 246 -4013 648 3947
rect 1068 3907 1868 3947
rect 1068 -3973 1468 3907
rect 1828 -3973 1868 3907
rect 1068 -4013 1868 -3973
rect 246 -4019 252 -4013
rect 206 -4031 252 -4019
<< via1 >>
rect -661 5317 -362 5616
rect 768 4867 1128 5227
rect -660 4338 -323 4675
rect -972 -3973 -612 3907
rect 1138 4337 1477 4676
rect 1468 -3973 1828 3907
<< metal2 >>
rect -661 5616 -362 5622
rect -1397 5322 -661 5612
rect -661 5311 -362 5317
rect 768 5227 1128 5233
rect 1128 4867 2228 5227
rect 768 4861 1128 4867
rect -660 4675 -323 4681
rect -1400 4338 -660 4675
rect -660 4332 -323 4338
rect 1138 4676 1477 4682
rect 1477 4337 2217 4676
rect 1138 4331 1477 4337
rect -1374 3907 -572 3947
rect -1374 -3973 -972 3907
rect -612 -3973 -572 3907
rect -1374 -4013 -572 -3973
rect 1426 3907 2228 3947
rect 1426 -3973 1468 3907
rect 1828 -3973 2228 3907
rect 1426 -4013 2228 -3973
<< labels >>
rlabel metal2 1828 -4013 2228 3947 3 D_Pin_L
<< properties >>
string FIXED_BBOX -363 -4162 363 4162
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 40 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
