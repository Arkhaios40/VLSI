* NGSPICE file created from AnalogFFT.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z a_n358_n1169# a_n492_n1391# a_n300_n1257#
+ a_300_n1169#
X0 a_300_n1169# a_n300_n1257# a_n358_n1169# a_n492_n1391# sky130_fd_pr__nfet_g5v0d10v5 ad=3.48e+12p pd=2.458e+07u as=3.48e+12p ps=2.458e+07u w=1.2e+07u l=3e+06u
.ends

.subckt NmosStage1 In Cp1 Cp2 GND
Xsky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_0 GND GND In In sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z
Xsky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_1 m1_n1260_n3620# GND In GND sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z
Xsky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_2 In GND In In sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z
Xsky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_3 Cp2 GND In m1_n1260_n3620# sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z
Xsky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_4 Cp1 GND In m1_n660_140# sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z
Xsky130_fd_pr__nfet_g5v0d10v5_CQJY2Z_5 m1_n660_140# GND In GND sky130_fd_pr__nfet_g5v0d10v5_CQJY2Z
C0 In GND 15.54fF
.ends

.subckt NMOSR2Stg1 Bit0i+ Out1 Bit0i- Out2 Out3 Out4 Out5 Bit1i- Out6 bit1q+ Out7
+ Bit1q- Out8 Bit0q- Bit1i+ VSUBS Bit0q+
XNmosStage1_0 Bit0i+ Out1 Out5 VSUBS NmosStage1
XNmosStage1_1 Bit1q- Out4 Out7 VSUBS NmosStage1
XNmosStage1_2 bit1q+ Out3 Out8 VSUBS NmosStage1
XNmosStage1_3 Bit1i- Out2 Out5 VSUBS NmosStage1
XNmosStage1_4 Bit1i+ Out1 Out6 VSUBS NmosStage1
XNmosStage1_5 Bit0q- Out4 Out8 VSUBS NmosStage1
XNmosStage1_6 Bit0q+ Out3 Out7 VSUBS NmosStage1
XNmosStage1_7 Bit0i- Out2 Out6 VSUBS NmosStage1
C0 Out5 Out7 10.23fF
C1 Out5 Out3 11.38fF
C2 Out8 Out7 25.76fF
C3 Out2 Out5 40.70fF
C4 Out8 Out5 10.28fF
C5 Out6 Out4 11.33fF
C6 Out6 Out7 10.56fF
C7 Out6 Out3 11.42fF
C8 Out6 Out5 20.73fF
C9 Out7 Out4 12.32fF
C10 Bit0i- VSUBS 13.65fF
C11 Bit0q+ VSUBS 13.53fF
C12 Bit0q- VSUBS 13.36fF
C13 Out1 VSUBS 39.92fF
C14 Out6 VSUBS 65.58fF
C15 Bit1i+ VSUBS 13.43fF
C16 Out2 VSUBS 43.23fF
C17 Out5 VSUBS 63.88fF
C18 Bit1i- VSUBS 13.64fF
C19 Out3 VSUBS 46.86fF
C20 Out8 VSUBS 80.92fF
C21 bit1q+ VSUBS 13.49fF
C22 Out4 VSUBS 50.88fF
C23 Out7 VSUBS 77.72fF
C24 Bit1q- VSUBS 13.59fF
C25 Bit0i+ VSUBS 13.77fF
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ a_n358_n1236# a_300_n1236# a_n300_n1262#
+ w_n558_n1462# VSUBS
X0 a_300_n1236# a_n300_n1262# a_n358_n1236# w_n558_n1462# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48e+12p pd=2.458e+07u as=3.48e+12p ps=2.458e+07u w=1.2e+07u l=3e+06u
C0 w_n558_n1462# VSUBS 10.98fF
.ends

.subckt Stage2Pmos In Cp2 Cp1 w_n2400_n180# VSUBS
Xsky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_0 In In In w_n2400_n180# VSUBS sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ
Xsky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_1 Cp2 m1_1408_2794# In w_n2400_n180# VSUBS sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ
Xsky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_2 w_n2400_n180# In In w_n2400_n180# VSUBS sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ
Xsky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_3 Cp1 m1_4640_2760# In w_n2400_n180# VSUBS sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ
Xsky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_4 m1_1408_2794# w_n2400_n180# In w_n2400_n180#
+ VSUBS sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ
Xsky130_fd_pr__pfet_g5v0d10v5_WNKUWZ_5 m1_4640_2760# w_n2400_n180# In w_n2400_n180#
+ VSUBS sky130_fd_pr__pfet_g5v0d10v5_WNKUWZ
C0 w_n2400_n180# In 16.67fF
C1 w_n2400_n180# VSUBS 135.64fF
.ends

.subckt PMOSOutStg In1 Y0_I+ In2 Y0_I- In3 Y0_Q+ In4 Y0_Q- In5 Y1_I+ In6 Y1_I- In7
+ Y1_Q+ In8 Y1_Q- In9 Y2_I+ In10 Y2_I- In11 Y2_Q+ In12 Y2_Q- Y3_I+ In14 Y3_I- In15
+ Y3_Q+ In16 Y3_Q- In13 VSUBS w_n2728_n8326#
XStage2Pmos_8 In8 Y3_Q- Y1_Q- w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_9 In7 Y3_Q+ Y1_Q+ w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_10 In1 Y2_I+ Y0_I+ w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_11 In5 Y3_I+ Y1_I+ w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_12 In4 Y2_Q- Y0_Q- w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_13 In3 Y2_Q+ Y0_Q+ w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_14 In2 Y2_I- Y0_I- w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_15 In16 Y3_Q+ Y1_Q- w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_0 In6 Y3_I- Y1_I- w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_1 In15 Y3_Q- Y1_Q+ w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_2 In14 Y3_I+ Y1_I- w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_3 In13 Y3_I- Y1_I+ w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_4 In12 Y2_Q+ Y0_Q- w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_5 In11 Y2_Q- Y0_Q+ w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_7 In9 Y2_I- Y0_I+ w_n2728_n8326# VSUBS Stage2Pmos
XStage2Pmos_6 In10 Y2_I+ Y0_I- w_n2728_n8326# VSUBS Stage2Pmos
C0 Y2_I- Y2_I+ 13.23fF
C1 Y0_I- VSUBS 52.81fF
C2 Y2_I+ VSUBS 40.03fF
C3 Y0_I+ VSUBS 50.64fF
C4 Y2_I- VSUBS 51.43fF
C5 Y0_Q+ VSUBS 52.57fF
C6 Y2_Q- VSUBS 57.78fF
C7 Y0_Q- VSUBS 54.30fF
C8 Y2_Q+ VSUBS 48.55fF
C9 In12 VSUBS 10.07fF
C10 Y1_I+ VSUBS 58.01fF
C11 Y3_I- VSUBS 62.17fF
C12 Y1_I- VSUBS 58.60fF
C13 Y3_I+ VSUBS 62.84fF
C14 Y1_Q+ VSUBS 60.74fF
C15 Y3_Q- VSUBS 69.82fF
C16 Y1_Q- VSUBS 62.71fF
C17 Y3_Q+ VSUBS 66.86fF
C18 w_n2728_n8326# VSUBS 725.83fF
.ends

.subckt AnalogFFT IN_X0_I+ OUT_Y0_I+ IN_X0_I- OUT_Y0_I- IN_X0_Q+ OUT_X0_Q+ IN_X0_Q-
+ OUT_X0_Q- IN_X2_I+ OUT_Y1_I+ IN_X2_I- OUT_Y1_I- IN_X2_Q+ OUT_Y1_Q+ IN_X2_Q- OUT_Y1_Q-
+ IN_X1_I+ OUT_Y2_I+ IN_X1_I- OUT_Y2_I- IN_X1_Q+ OUT_Y2_Q+ IN_X1_Q- OUT_Y2_Q- IN_X3_I+
+ OUT_Y3_I+ IN_X3_I- OUT_Y3_I- IN_X3_Q+ OUT_Y3_Q+ IN_X3_Q- OUT_Y3_Q-
XNMOSR2Stg1_1 IN_X1_I+ PMOSOutStg_0/In9 IN_X1_I- PMOSOutStg_0/In10 PMOSOutStg_0/In11
+ PMOSOutStg_0/In12 PMOSOutStg_0/In13 IN_X3_I- PMOSOutStg_0/In14 IN_X3_Q+ PMOSOutStg_0/In15
+ IN_X3_Q- PMOSOutStg_0/In16 IN_X1_Q- IN_X3_I+ GND IN_X1_Q+ NMOSR2Stg1
XPMOSOutStg_0 PMOSOutStg_0/In1 OUT_Y0_I+ PMOSOutStg_0/In2 OUT_Y0_I- PMOSOutStg_0/In3
+ OUT_X0_Q+ PMOSOutStg_0/In4 OUT_X0_Q- PMOSOutStg_0/In5 OUT_Y1_I+ PMOSOutStg_0/In6
+ OUT_Y1_I- PMOSOutStg_0/In7 OUT_Y1_Q+ PMOSOutStg_0/In8 OUT_Y1_Q- PMOSOutStg_0/In9
+ OUT_Y2_I+ PMOSOutStg_0/In10 OUT_Y2_I- PMOSOutStg_0/In11 OUT_Y2_Q+ PMOSOutStg_0/In12
+ OUT_Y2_Q- OUT_Y3_I+ PMOSOutStg_0/In14 OUT_Y3_I- PMOSOutStg_0/In15 OUT_Y3_Q+ PMOSOutStg_0/In16
+ OUT_Y3_Q- PMOSOutStg_0/In13 GND Vdd PMOSOutStg
XNMOSR2Stg1_0 IN_X0_I+ PMOSOutStg_0/In1 IN_X0_I- PMOSOutStg_0/In2 PMOSOutStg_0/In3
+ PMOSOutStg_0/In4 PMOSOutStg_0/In5 IN_X2_I- PMOSOutStg_0/In6 IN_X2_Q+ PMOSOutStg_0/In7
+ IN_X2_Q- PMOSOutStg_0/In8 IN_X0_Q- IN_X2_I+ GND IN_X0_Q+ NMOSR2Stg1
C0 IN_X0_I- GND 21.08fF
C1 IN_X0_Q+ GND 20.87fF
C2 IN_X0_Q- GND 20.69fF
C3 IN_X2_I+ GND 20.74fF
C4 IN_X2_I- GND 20.90fF
C5 IN_X2_Q+ GND 20.57fF
C6 IN_X2_Q- GND 20.62fF
C7 IN_X0_I+ GND 17.69fF
C8 OUT_Y0_I- GND 58.72fF
C9 OUT_Y2_I+ GND 51.02fF
C10 PMOSOutStg_0/In10 GND 81.88fF
C11 OUT_Y0_I+ GND 57.67fF
C12 OUT_Y2_I- GND 59.48fF
C13 PMOSOutStg_0/In9 GND 81.71fF
C14 OUT_X0_Q+ GND 58.50fF
C15 OUT_Y2_Q- GND 66.92fF
C16 PMOSOutStg_0/In11 GND 85.43fF
C17 OUT_X0_Q- GND 60.28fF
C18 OUT_Y2_Q+ GND 57.60fF
C19 PMOSOutStg_0/In12 GND 88.38fF
C20 OUT_Y1_I+ GND 64.27fF
C21 OUT_Y3_I- GND 70.63fF
C22 PMOSOutStg_0/In13 GND 110.60fF
C23 OUT_Y1_I- GND 63.85fF
C24 OUT_Y3_I+ GND 73.24fF
C25 PMOSOutStg_0/In14 GND 111.63fF
C26 OUT_Y1_Q+ GND 66.10fF
C27 OUT_Y3_Q- GND 77.42fF
C28 PMOSOutStg_0/In15 GND 123.62fF
C29 PMOSOutStg_0/In6 GND 103.52fF
C30 OUT_Y1_Q- GND 68.30fF
C31 OUT_Y3_Q+ GND 74.95fF
C32 PMOSOutStg_0/In16 GND 121.63fF
C33 Vdd GND -457.86fF
C34 PMOSOutStg_0/In2 GND 86.34fF
C35 PMOSOutStg_0/In3 GND 92.38fF
C36 PMOSOutStg_0/In4 GND 96.06fF
C37 PMOSOutStg_0/In5 GND 102.19fF
C38 PMOSOutStg_0/In1 GND 74.50fF
C39 PMOSOutStg_0/In7 GND 116.13fF
C40 PMOSOutStg_0/In8 GND 119.96fF
C41 IN_X1_I- GND 21.56fF
C42 IN_X1_Q+ GND 20.90fF
C43 IN_X1_Q- GND 20.69fF
C44 IN_X3_I+ GND 20.74fF
C45 IN_X3_I- GND 20.88fF
C46 IN_X3_Q+ GND 20.58fF
C47 IN_X3_Q- GND 20.61fF
C48 IN_X1_I+ GND 21.38fF
.ends

