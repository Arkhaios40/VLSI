* NGSPICE file created from OpAmp.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_g5v0d10v5_97BMAW a_n558_n3000# a_n500_n3097# a_500_n3000#
+ w_n758_n3297#
X0 a_500_n3000# a_n500_n3097# a_n558_n3000# w_n758_n3297# sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+12p pd=6.058e+07u as=8.7e+12p ps=6.058e+07u w=3e+07u l=5e+06u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_97TZA6 a_n200_n2097# a_200_n2000# w_n458_n2297#
+ a_n258_n2000#
X0 a_200_n2000# a_n200_n2097# a_n258_n2000# w_n458_n2297# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=2e+06u
.ends

.subckt PMOSPair body CenterTap Vp m1_162_3398# Vs
XXM12 Vs Vp CenterTap body sky130_fd_pr__pfet_g5v0d10v5_97BMAW
XXM7 Vp CenterTap body m1_162_3398# sky130_fd_pr__pfet_g5v0d10v5_97TZA6
XXM8 Vp m1_162_3398# body CenterTap sky130_fd_pr__pfet_g5v0d10v5_97TZA6
XXM9 Vp CenterTap body m1_162_3398# sky130_fd_pr__pfet_g5v0d10v5_97TZA6
XXM10 Vp m1_162_3398# body CenterTap sky130_fd_pr__pfet_g5v0d10v5_97TZA6
XXM11 Vp CenterTap body m1_162_3398# sky130_fd_pr__pfet_g5v0d10v5_97TZA6
.ends

.subckt ConnectedPMOSPair Vss VP_LeftPin R_Pin
XPMOSPair_0 Vss PMOSPair_0/CenterTap VP_LeftPin R_Pin Vss PMOSPair
XPMOSPair_1 Vss PMOSPair_1/CenterTap VP_LeftPin VP_LeftPin Vss PMOSPair
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UBJTTH D_Pin_L a_n258_n4031# li_688_4007# a_n392_n4191#
+ a_n200_n4057# a_200_n4031#
X0 a_200_n4031# a_n200_n4057# a_n258_n4031# a_n392_n4191# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16e+13p pd=8.058e+07u as=1.16e+13p ps=8.058e+07u w=4e+07u l=2e+06u
.ends

.subckt DifferentialPair D_Pin_R D_In_L D_In_R NMOS_Vs Body D_Pin_L
Xsky130_fd_pr__nfet_g5v0d10v5_UBJTTH_0 D_Pin_L D_Pin_R D_In_L Body D_In_R NMOS_Vs
+ sky130_fd_pr__nfet_g5v0d10v5_UBJTTH
X0 NMOS_Vs D_In_L D_Pin_L Body sky130_fd_pr__nfet_g5v0d10v5 ad=2.28172e+13p pd=1.58815e+08u as=1.16e+13p ps=8.058e+07u w=4e+07u l=2e+06u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2ZQVB2 a_n492_n2191# li_n480_2135# a_n300_n2057#
+ a_300_n2031# a_n358_n2031#
X0 a_300_n2031# a_n300_n2057# a_n358_n2031# a_n492_n2191# sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=3e+06u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_49CJ6G a_n108_n2531# a_n242_n2691# a_50_n2531#
+ a_n50_n2557#
X0 a_50_n2531# a_n50_n2557# a_n108_n2531# a_n242_n2691# sky130_fd_pr__nfet_g5v0d10v5 ad=7.25e+12p pd=5.058e+07u as=7.25e+12p ps=5.058e+07u w=2.5e+07u l=500000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_M768YF li_n398_3150# a_500_n3036# a_n500_n3062#
+ w_n758_n3262# a_n558_n3036#
X0 a_500_n3036# a_n500_n3062# a_n558_n3036# w_n758_n3262# sky130_fd_pr__pfet_g5v0d10v5 ad=8.7e+12p pd=6.058e+07u as=8.7e+12p ps=6.058e+07u w=3e+07u l=5e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_27X89E m3_n1186_n540# c1_n1146_n500#
X0 c1_n1146_n500# m3_n1186_n540# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=1e+07u
.ends

.subckt GainStage VPlus Gain_L_Pin Gain_R_Pin GateRef Out Gain_Vs
Xsky130_fd_pr__nfet_g5v0d10v5_2ZQVB2_1 Gain_Vs Gain_L_Pin Gain_L_Pin Gain_Vs Gain_L_Pin
+ sky130_fd_pr__nfet_g5v0d10v5_2ZQVB2
Xsky130_fd_pr__nfet_g5v0d10v5_49CJ6G_0 Gain_Vs Gain_Vs Out Gain_R_Pin sky130_fd_pr__nfet_g5v0d10v5_49CJ6G
Xsky130_fd_pr__nfet_g5v0d10v5_49CJ6G_1 Out Gain_Vs Gain_Vs Gain_R_Pin sky130_fd_pr__nfet_g5v0d10v5_49CJ6G
Xsky130_fd_pr__pfet_g5v0d10v5_M768YF_0 GateRef VPlus GateRef VPlus Out sky130_fd_pr__pfet_g5v0d10v5_M768YF
Xsky130_fd_pr__pfet_g5v0d10v5_M768YF_1 GateRef Out GateRef VPlus VPlus sky130_fd_pr__pfet_g5v0d10v5_M768YF
Xsky130_fd_pr__pfet_g5v0d10v5_M768YF_2 GateRef VPlus GateRef VPlus Out sky130_fd_pr__pfet_g5v0d10v5_M768YF
Xsky130_fd_pr__cap_mim_m3_1_27X89E_0 Gain_R_Pin Out sky130_fd_pr__cap_mim_m3_1
Xsky130_fd_pr__nfet_g5v0d10v5_2ZQVB2_0 Gain_Vs Gain_Vs Gain_L_Pin Gain_R_Pin Gain_Vs
+ sky130_fd_pr__nfet_g5v0d10v5_2ZQVB2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HYQESV a_200_n2031# a_n258_n2031# a_n392_n2191#
+ a_n200_n2057#
X0 a_200_n2031# a_n200_n2057# a_n258_n2031# a_n392_n2191# sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+12p pd=4.058e+07u as=5.8e+12p ps=4.058e+07u w=2e+07u l=2e+06u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_VSVLYK a_n558_n1031# a_n692_n1191# a_n500_n1057#
+ a_500_n1031#
X0 a_500_n1031# a_n500_n1057# a_n558_n1031# a_n692_n1191# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p ps=2.058e+07u w=1e+07u l=5e+06u
.ends

.subckt NMOSPair Vd Vn S VSUBS
Xsky130_fd_pr__nfet_g5v0d10v5_HYQESV_0 m1_n2132_2872# Vd VSUBS Vn sky130_fd_pr__nfet_g5v0d10v5_HYQESV
Xsky130_fd_pr__nfet_g5v0d10v5_HYQESV_1 m1_n2132_2872# Vd VSUBS Vn sky130_fd_pr__nfet_g5v0d10v5_HYQESV
Xsky130_fd_pr__nfet_g5v0d10v5_VSVLYK_0 S VSUBS Vn Vd sky130_fd_pr__nfet_g5v0d10v5_VSVLYK
Xsky130_fd_pr__nfet_g5v0d10v5_HYQESV_2 Vd m1_n2132_2872# VSUBS Vn sky130_fd_pr__nfet_g5v0d10v5_HYQESV
Xsky130_fd_pr__nfet_g5v0d10v5_HYQESV_3 m1_n2132_2872# Vd VSUBS Vn sky130_fd_pr__nfet_g5v0d10v5_HYQESV
Xsky130_fd_pr__nfet_g5v0d10v5_HYQESV_4 Vd m1_n2132_2872# VSUBS Vn sky130_fd_pr__nfet_g5v0d10v5_HYQESV
.ends

.subckt ConnectedNMOSPair R_Pin L_Pin Vs
XNMOSPair_0 R_Pin L_Pin Vs Vs NMOSPair
XNMOSPair_1 L_Pin L_Pin Vs Vs NMOSPair
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_3ZBBQK a_n3862_n4398# a_3450_n4268# a_n3732_n4268#
X0 a_n3732_n4268# a_3450_n4268# a_n3862_n4398# sky130_fd_pr__res_xhigh_po w=1.41e+06u l=7.8337e+08u
.ends

.subckt CurRefResistor Pin1 Pin2
Xsky130_fd_pr__res_xhigh_po_1p41_3ZBBQK_0 VSUBS Pin2 Pin1 sky130_fd_pr__res_xhigh_po_1p41
.ends

.subckt CurrentRef Vplus Ref Vneg
XCurRefResistor_0 Vplus CurRefResistor_0/Pin2 CurRefResistor
XConnectedNMOSPair_0 Ref CurRefResistor_0/Pin2 Vneg ConnectedNMOSPair
.ends

*.subckt OpAmp VDD In+ In- Out Ground
XConnectedPMOSPair_1 VDD PMOSPair_1/Vp ConnectedPMOSPair_1/R_Pin ConnectedPMOSPair
XPMOSPair_0 VDD PMOSPair_0/CenterTap PMOSPair_1/Vp GainStage_0/Gain_L_Pin VDD PMOSPair
XPMOSPair_1 VDD PMOSPair_1/CenterTap PMOSPair_1/Vp GainStage_0/Gain_R_Pin VDD PMOSPair
XDifferentialPair_0 PMOSPair_1/CenterTap In+ In- ConnectedNMOSPair_0/R_Pin Ground
+ PMOSPair_0/CenterTap DifferentialPair
XGainStage_0 VDD GainStage_0/Gain_L_Pin GainStage_0/Gain_R_Pin PMOSPair_1/Vp Out Ground
+ GainStage
XConnectedNMOSPair_0 ConnectedNMOSPair_0/R_Pin ConnectedPMOSPair_1/R_Pin Ground ConnectedNMOSPair
XCurrentRef_0 VDD PMOSPair_1/Vp Ground CurrentRef
*.ends

