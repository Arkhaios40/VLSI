magic
tech sky130A
magscale 1 2
timestamp 1670438645
<< nwell >>
rect -2714 -1938 10852 89584
rect -2728 -8326 10902 -1938
<< viali >>
rect 25251 77067 25905 77721
<< metal1 >>
rect 8050 85240 10976 85276
rect 6340 85141 10976 85240
rect 6340 84487 9729 85141
rect 10383 85092 10976 85141
rect 10383 84487 35715 85092
rect 6340 84438 35715 84487
rect 6340 84374 10976 84438
rect 6340 84302 10554 84374
rect -5684 83086 1318 84234
rect 3560 83905 10554 84006
rect 35061 83911 35715 84438
rect 20675 83905 21329 83911
rect 3560 83251 20675 83905
rect 3560 83050 10554 83251
rect 20675 83245 21329 83251
rect 35059 83905 35715 83911
rect 35713 83251 35715 83905
rect 35059 83245 35715 83251
rect 35061 83239 35715 83245
rect 6432 79217 10646 79406
rect 6432 78552 13065 79217
rect 13730 78552 35672 79217
rect 6432 78468 10646 78552
rect -5822 77230 1958 78378
rect 3652 77721 10646 78062
rect 25206 77721 26010 77794
rect 35007 77727 35672 78552
rect 3652 77106 25251 77721
rect 9671 77067 25251 77106
rect 25905 77067 26010 77721
rect 25206 76942 26010 77067
rect 34897 77721 35672 77727
rect 35551 77268 35672 77721
rect 34897 77061 35551 77067
rect 6432 73408 10646 73590
rect 6432 72710 14329 73408
rect 15027 72710 35881 73408
rect 6432 72652 10646 72710
rect -5794 71354 1986 72502
rect 3652 72179 10646 72338
rect 35183 72185 35881 72710
rect 26457 72179 27111 72185
rect 3652 71525 26457 72179
rect 3652 71382 10646 71525
rect 26457 71519 27111 71525
rect 35059 72179 35881 72185
rect 35713 71525 35881 72179
rect 35059 71519 35881 71525
rect 35183 71379 35881 71519
rect 6468 67491 10682 67700
rect 6468 66865 15519 67491
rect 16145 66865 31357 67491
rect -5878 65618 1902 66766
rect 6468 66762 10682 66865
rect 3670 66315 10664 66466
rect 30731 66412 31357 66865
rect 27661 66315 28315 66321
rect 3670 65661 27661 66315
rect 3670 65510 10664 65661
rect 27661 65655 28315 65661
rect 30566 66315 31486 66412
rect 30566 65661 30597 66315
rect 31251 65661 31486 66315
rect 30566 65604 31486 65661
rect 6266 61522 10480 61682
rect 6266 60868 17197 61522
rect 17851 60868 35401 61522
rect 6266 60744 10480 60868
rect -6076 59518 1704 60666
rect 3524 60213 10518 60412
rect 29188 60213 30094 60358
rect 34747 60219 35401 60868
rect 3524 59559 29267 60213
rect 29921 59559 30094 60213
rect 3524 59456 10518 59559
rect 29188 59432 30094 59559
rect 34735 60213 35401 60219
rect 35389 59559 35401 60213
rect 34735 59553 35401 59559
rect 34747 59539 35401 59553
rect 6302 55132 10516 55334
rect 6302 54506 18603 55132
rect 19229 54506 35221 55132
rect 6302 54396 10516 54506
rect -6076 53164 1704 54312
rect 9698 54062 10324 54064
rect 3504 53707 10498 54062
rect 34595 53964 35221 54506
rect 30578 53707 31484 53854
rect 3504 53106 30713 53707
rect 9671 53053 30713 53106
rect 31367 53053 31484 53707
rect 30578 52928 31484 53053
rect 34500 53707 35500 53964
rect 34500 53053 34653 53707
rect 35307 53053 35500 53707
rect 34500 52796 35500 53053
rect 6376 49530 10590 49664
rect 19890 49530 20890 49654
rect 6376 48876 20021 49530
rect 20675 48876 35345 49530
rect 6376 48726 10590 48876
rect 19890 48760 20890 48876
rect -6048 47512 1732 48660
rect 3596 48165 10590 48450
rect 32046 48165 32952 48256
rect 3596 47511 32159 48165
rect 32813 47511 32952 48165
rect 34691 48171 35345 48876
rect 34691 48165 35389 48171
rect 34691 47515 34735 48165
rect 3596 47494 10590 47511
rect 32046 47330 32952 47511
rect 34735 47505 35389 47511
rect 6412 43546 10626 43830
rect 21410 43546 22558 43776
rect 34505 43546 35131 43552
rect 6412 42920 21763 43546
rect 22389 42920 34505 43546
rect 6412 42892 10626 42920
rect -6048 41692 1732 42840
rect 21410 42782 22558 42920
rect 34505 42914 35131 42920
rect 3634 42289 10628 42542
rect 21578 42289 22232 42296
rect 33699 42289 34325 42295
rect 3634 41663 33699 42289
rect 3634 41586 10628 41663
rect 21578 40302 22232 41663
rect 33699 41657 34325 41663
rect 6486 37598 10700 37794
rect 6486 36936 9766 37598
rect 10428 36936 10700 37598
rect 6486 36856 10700 36936
rect -6076 35592 1704 36740
rect 3616 36370 10610 36506
rect 3616 35716 9783 36370
rect 10437 35716 10610 36370
rect 3616 35550 10610 35716
rect 6596 31372 10810 31482
rect 6596 30712 9736 31372
rect 10396 30712 10810 31372
rect 6596 30544 10810 30712
rect -5992 29378 1788 30526
rect 9780 30248 10674 30288
rect 3726 30156 10720 30248
rect 3726 29502 9910 30156
rect 10564 29502 10720 30156
rect 3726 29292 10720 29502
rect 6524 25296 10738 25446
rect 6524 24642 9885 25296
rect 10539 24642 10738 25296
rect 6524 24508 10738 24642
rect -6104 23278 1676 24426
rect 3726 24074 10720 24174
rect 3726 23420 12555 24074
rect 3726 23218 10720 23420
rect 6468 19176 10682 19336
rect 6468 18522 9727 19176
rect 10381 18522 10682 19176
rect 6468 18398 10682 18522
rect -6188 17176 1592 18324
rect 3634 17954 10628 18102
rect 3634 17300 9826 17954
rect 10480 17300 10628 17954
rect 11901 17961 12555 23420
rect 15353 17961 16007 17967
rect 11901 17307 15353 17961
rect 15353 17301 16007 17307
rect 3634 17146 10628 17300
rect 9708 17128 10602 17146
rect 6486 13492 10700 13666
rect 6486 12838 9898 13492
rect 10552 12838 10700 13492
rect 6486 12728 10700 12838
rect -5878 11470 1902 12618
rect 3762 12270 10756 12342
rect 14060 12270 14900 12354
rect 3762 11616 14123 12270
rect 14777 11616 14900 12270
rect 3762 11386 10756 11616
rect 14060 11502 14900 11616
rect 15792 12239 16632 12334
rect 15792 11585 15881 12239
rect 16535 11585 16632 12239
rect 15792 11482 16632 11585
rect 15881 9935 16535 11482
rect 12521 9281 16535 9935
rect 6578 7676 10792 7796
rect 6578 7022 10060 7676
rect 10714 7022 10792 7676
rect 6578 6858 10792 7022
rect -5794 5622 1986 6770
rect 3910 6454 10904 6654
rect 12521 6454 13175 9281
rect 3910 5800 13175 6454
rect 3910 5698 10904 5800
rect 6652 2318 10866 2514
rect 6652 1664 10105 2318
rect 10759 1664 10866 2318
rect 6652 1576 10866 1664
rect -5682 252 2098 1400
rect 3946 1133 10940 1208
rect 13941 1133 14567 1139
rect 3946 507 13941 1133
rect 3946 252 10940 507
rect 13941 501 14567 507
rect 16383 377 16389 1031
rect 17043 377 17049 1031
rect 6854 -3926 11088 -3780
rect 6854 -4580 10212 -3926
rect 10866 -4580 11088 -3926
rect 6854 -4682 11088 -4580
rect -5514 -5934 2266 -4786
rect 4038 -5148 11032 -5032
rect 16389 -5148 17043 377
rect 4038 -5802 17043 -5148
rect 4038 -5988 11032 -5802
<< via1 >>
rect 9729 84487 10383 85141
rect 20675 83251 21329 83905
rect 35059 83251 35713 83905
rect 13065 78552 13730 79217
rect 25251 77067 25905 77721
rect 34897 77067 35551 77721
rect 14329 72710 15027 73408
rect 26457 71525 27111 72179
rect 35059 71525 35713 72179
rect 15519 66865 16145 67491
rect 27661 65661 28315 66315
rect 30597 65661 31251 66315
rect 17197 60868 17851 61522
rect 29267 59559 29921 60213
rect 34735 59559 35389 60213
rect 18603 54506 19229 55132
rect 30713 53053 31367 53707
rect 34653 53053 35307 53707
rect 20021 48876 20675 49530
rect 32159 47511 32813 48165
rect 34735 47511 35389 48165
rect 21763 42920 22389 43546
rect 34505 42920 35131 43546
rect 33699 41663 34325 42289
rect 9766 36936 10428 37598
rect 9783 35716 10437 36370
rect 9736 30712 10396 31372
rect 9910 29502 10564 30156
rect 9885 24642 10539 25296
rect 9727 18522 10381 19176
rect 9826 17300 10480 17954
rect 15353 17307 16007 17961
rect 9898 12838 10552 13492
rect 14123 11616 14777 12270
rect 15881 11585 16535 12239
rect 10060 7022 10714 7676
rect 10105 1664 10759 2318
rect 13941 507 14567 1133
rect 16389 377 17043 1031
rect 10212 -4580 10866 -3926
<< metal2 >>
rect 9729 85141 10383 85147
rect 11624 85141 12278 85142
rect 10383 84487 12278 85141
rect 9729 84481 10383 84487
rect 9692 37598 10458 37632
rect 9692 36936 9766 37598
rect 10428 37596 10458 37598
rect 11624 37596 12278 84487
rect 23908 83905 24552 83909
rect 20669 83251 20675 83905
rect 21329 83900 24557 83905
rect 21329 83256 23908 83900
rect 24552 83256 24557 83900
rect 21329 83251 24557 83256
rect 35053 83251 35059 83905
rect 35713 83251 36681 83905
rect 37335 83251 37344 83905
rect 23908 83247 24552 83251
rect 13065 79217 13730 79223
rect 13039 78552 13065 79057
rect 13039 78546 13730 78552
rect 10428 36939 12280 37596
rect 10428 36936 10458 36939
rect 9692 36862 10458 36936
rect 9783 36370 10437 36376
rect 9774 35716 9783 36370
rect 10437 35716 10446 36370
rect 9783 35710 10437 35716
rect 9672 31372 10584 31414
rect 9672 30712 9736 31372
rect 10396 31370 10584 31372
rect 13039 31370 13693 78546
rect 25206 77721 26010 77794
rect 25206 77067 25251 77721
rect 25905 77067 26010 77721
rect 34891 77067 34897 77721
rect 35551 77067 36681 77721
rect 37335 77067 37344 77721
rect 25206 76942 26010 77067
rect 14329 73408 15027 73414
rect 14329 72704 15027 72710
rect 10396 30714 13694 31370
rect 10396 30712 10584 30714
rect 9672 30664 10584 30712
rect 9780 30156 10674 30288
rect 9780 29502 9910 30156
rect 10564 29502 10674 30156
rect 9780 29344 10674 29502
rect 9885 25296 10539 25302
rect 14336 25296 14992 72704
rect 26462 72179 27106 72183
rect 26451 71525 26457 72179
rect 27111 71525 27117 72179
rect 35053 71525 35059 72179
rect 35713 71525 36033 72179
rect 36687 71525 36696 72179
rect 26462 71521 27106 71525
rect 10539 24642 14992 25296
rect 9885 24636 10539 24642
rect 14336 24641 14992 24642
rect 15427 67497 16081 67701
rect 15427 67491 16145 67497
rect 15427 66865 15519 67491
rect 15427 66859 16145 66865
rect 9616 19176 10490 19318
rect 15427 19176 16081 66859
rect 27666 66315 28310 66319
rect 30566 66315 31486 66412
rect 35789 66315 36443 66324
rect 27655 65661 27661 66315
rect 28315 65661 28321 66315
rect 30566 65661 30597 66315
rect 31251 65661 35789 66315
rect 27666 65657 28310 65661
rect 30566 65604 31486 65661
rect 35789 65652 36443 65661
rect 17235 61528 17889 61623
rect 17197 61522 17889 61528
rect 17851 60868 17889 61522
rect 17197 60862 17889 60868
rect 9616 18522 9727 19176
rect 10381 18522 16169 19176
rect 9616 18408 10490 18522
rect 9708 17954 10602 18072
rect 9708 17300 9826 17954
rect 10480 17300 10602 17954
rect 9708 17128 10602 17300
rect 15222 17961 16116 18112
rect 15222 17307 15353 17961
rect 16007 17307 16116 17961
rect 15222 17168 16116 17307
rect 9820 13492 10656 13584
rect 17235 13492 17889 60862
rect 29188 60213 30094 60358
rect 29188 59559 29267 60213
rect 29921 59559 30094 60213
rect 34729 59559 34735 60213
rect 35389 59559 35869 60213
rect 36523 59559 36532 60213
rect 29188 59432 30094 59559
rect 9820 12838 9898 13492
rect 10552 12838 17889 13492
rect 18569 55138 19223 55421
rect 18569 55132 19229 55138
rect 18569 54506 18603 55132
rect 18569 54500 19229 54506
rect 9820 12716 10656 12838
rect 14060 12270 14900 12354
rect 14060 11616 14123 12270
rect 14777 11616 14900 12270
rect 14060 11502 14900 11616
rect 15792 12239 16632 12334
rect 15792 11585 15881 12239
rect 16535 11585 16632 12239
rect 15792 11482 16632 11585
rect 9988 7676 10720 7740
rect 18569 7676 19223 54500
rect 30578 53707 31484 53854
rect 30578 53053 30713 53707
rect 31367 53053 31484 53707
rect 30578 52928 31484 53053
rect 34653 53707 35307 53713
rect 35307 53053 36195 53707
rect 36849 53053 36858 53707
rect 34653 53047 35307 53053
rect 19890 49530 20890 49654
rect 19890 48876 20021 49530
rect 20675 48876 20890 49530
rect 19890 48760 20890 48876
rect 9988 7022 10060 7676
rect 10714 7022 19223 7676
rect 9988 6924 10720 7022
rect 10030 2318 10762 2408
rect 20069 2318 20723 48760
rect 32046 48165 32952 48256
rect 32046 47511 32159 48165
rect 32813 47511 32952 48165
rect 34729 47511 34735 48165
rect 35389 47511 36195 48165
rect 36849 47511 36858 48165
rect 32046 47330 32952 47511
rect 21568 43546 22450 43694
rect 21568 42920 21763 43546
rect 22389 42920 22450 43546
rect 34496 42920 34505 43546
rect 35131 42920 35140 43546
rect 21568 42802 22450 42920
rect 10030 1664 10105 2318
rect 10759 1664 20723 2318
rect 10030 1592 10762 1664
rect 13941 1133 14567 1142
rect 13935 507 13941 1133
rect 14567 507 14573 1133
rect 16389 1031 17043 1037
rect 13941 498 14567 507
rect 16380 377 16389 1031
rect 17043 377 17052 1031
rect 16389 371 17043 377
rect 10124 -3926 10856 -3832
rect 21653 -3926 22307 42802
rect 33704 42289 34320 42293
rect 33693 41663 33699 42289
rect 34325 41663 34331 42289
rect 33704 41659 34320 41663
rect 10124 -4580 10212 -3926
rect 10866 -4580 22307 -3926
rect 10124 -4648 10856 -4580
<< via2 >>
rect 23908 83256 24552 83900
rect 36681 83251 37335 83905
rect 9783 35716 10437 36370
rect 25256 77072 25900 77716
rect 36681 77067 37335 77721
rect 9910 29502 10564 30156
rect 26462 71530 27106 72174
rect 36033 71525 36687 72179
rect 27666 65666 28310 66310
rect 35789 65661 36443 66315
rect 9826 17300 10480 17954
rect 15353 17307 16007 17961
rect 29272 59564 29916 60208
rect 35869 59559 36523 60213
rect 14123 11616 14777 12270
rect 15881 11585 16535 12239
rect 30718 53058 31362 53702
rect 36195 53053 36849 53707
rect 32164 47516 32808 48160
rect 36195 47511 36849 48165
rect 34505 42920 35131 43546
rect 13941 507 14567 1133
rect 16389 377 17043 1031
rect 33704 41668 34320 42284
<< metal3 >>
rect 23904 83905 24556 83910
rect 36676 83905 37340 83910
rect 40087 83905 40741 83911
rect 23903 83904 24557 83905
rect 23903 83252 23904 83904
rect 24556 83252 24557 83904
rect 23903 83251 24557 83252
rect 36676 83251 36681 83905
rect 37335 83251 40087 83905
rect 23904 83246 24556 83251
rect 36676 83246 37340 83251
rect 40087 83245 40741 83251
rect 25206 77716 26010 77794
rect 25206 77072 25256 77716
rect 25900 77072 26010 77716
rect 25206 76942 26010 77072
rect 36676 77721 37340 77726
rect 39925 77721 40579 77727
rect 36676 77067 36681 77721
rect 37335 77067 39925 77721
rect 36676 77062 37340 77067
rect 39925 77061 40579 77067
rect 9778 36370 10442 36375
rect 9778 35716 9783 36370
rect 10437 35716 12281 36370
rect 9778 35711 10442 35716
rect 9780 30161 10674 30288
rect 9780 29497 9905 30161
rect 10569 29497 10674 30161
rect 9780 29344 10674 29497
rect 11627 30119 12281 35716
rect 25251 30286 25905 76942
rect 36028 72179 36692 72184
rect 39763 72179 40417 72185
rect 26457 72174 27111 72179
rect 26457 71530 26462 72174
rect 27106 71530 27111 72174
rect 25150 30119 26004 30286
rect 11627 29465 25251 30119
rect 25905 29465 26004 30119
rect 25150 29286 26004 29465
rect 26457 24079 27111 71530
rect 36028 71525 36033 72179
rect 36687 71525 39763 72179
rect 36028 71520 36692 71525
rect 39763 71519 40417 71525
rect 35784 66315 36448 66320
rect 13275 23425 26381 24079
rect 27035 23425 27111 24079
rect 27661 66310 28315 66315
rect 27661 65666 27666 66310
rect 28310 65666 28315 66310
rect 9708 17954 10602 18072
rect 13275 17954 13929 23425
rect 9708 17300 9826 17954
rect 10480 17300 13929 17954
rect 15222 17961 16116 18112
rect 27661 17961 28315 65666
rect 35784 65661 35789 66315
rect 36443 65661 39683 66315
rect 40337 65661 40343 66315
rect 35784 65656 36448 65661
rect 29267 60358 29921 60373
rect 29188 60208 30094 60358
rect 29188 59564 29272 60208
rect 29916 59564 30094 60208
rect 29188 59432 30094 59564
rect 35864 60213 36528 60218
rect 35864 59559 35869 60213
rect 36523 59559 39763 60213
rect 40417 59559 40423 60213
rect 35864 59554 36528 59559
rect 15222 17307 15353 17961
rect 16007 17307 27515 17961
rect 28169 17307 28315 17961
rect 9708 17128 10602 17300
rect 15222 17168 16116 17307
rect 14118 12270 14782 12275
rect 14118 11616 14123 12270
rect 14777 11616 14782 12270
rect 14118 11611 14782 11616
rect 15792 12239 16632 12334
rect 29267 12239 29921 59432
rect 30578 53702 31484 53854
rect 30578 53058 30718 53702
rect 31362 53058 31484 53702
rect 30578 52928 31484 53058
rect 36190 53707 36854 53712
rect 36190 53053 36195 53707
rect 36849 53053 39763 53707
rect 40417 53053 40423 53707
rect 36190 53048 36854 53053
rect 14123 6341 14777 11611
rect 15792 11585 15881 12239
rect 16535 11585 29057 12239
rect 29711 11585 29921 12239
rect 15792 11482 16632 11585
rect 30713 6508 31367 52928
rect 32046 48160 32952 48256
rect 32046 47516 32164 48160
rect 32808 47516 32952 48160
rect 32046 47330 32952 47516
rect 36190 48165 36854 48170
rect 36190 47511 36195 48165
rect 36849 47511 39519 48165
rect 40173 47511 40179 48165
rect 36190 47506 36854 47511
rect 30318 6341 31367 6508
rect 14123 5687 30435 6341
rect 31089 5687 31367 6341
rect 30318 5550 31226 5687
rect 32159 1180 32813 47330
rect 34500 43546 35136 43551
rect 34500 42920 34505 43546
rect 35131 42920 41805 43546
rect 42431 42920 42437 43546
rect 34500 42915 35136 42920
rect 13936 1133 14572 1138
rect 13936 507 13941 1133
rect 14567 507 14572 1133
rect 13936 502 14572 507
rect 16384 1031 17048 1036
rect 31884 1031 32813 1180
rect 13941 -1639 14567 502
rect 16384 377 16389 1031
rect 17043 377 31977 1031
rect 32631 377 32813 1031
rect 33699 42284 34325 42289
rect 33699 41668 33704 42284
rect 34320 41668 34325 42284
rect 16384 372 17048 377
rect 31884 222 32792 377
rect 13941 -2265 19645 -1639
rect 19019 -5389 19645 -2265
rect 33699 -5282 34325 41668
rect 33574 -5389 34450 -5282
rect 19019 -6015 33699 -5389
rect 34325 -6015 34450 -5389
rect 33574 -6138 34450 -6015
<< via3 >>
rect 23904 83900 24556 83904
rect 23904 83256 23908 83900
rect 23908 83256 24552 83900
rect 24552 83256 24556 83900
rect 23904 83252 24556 83256
rect 40087 83251 40741 83905
rect 39925 77067 40579 77721
rect 9905 30156 10569 30161
rect 9905 29502 9910 30156
rect 9910 29502 10564 30156
rect 10564 29502 10569 30156
rect 9905 29497 10569 29502
rect 25251 29465 25905 30119
rect 39763 71525 40417 72179
rect 26381 23425 27035 24079
rect 39683 65661 40337 66315
rect 39763 59559 40417 60213
rect 27515 17307 28169 17961
rect 39763 53053 40417 53707
rect 29057 11585 29711 12239
rect 39519 47511 40173 48165
rect 30435 5687 31089 6341
rect 41805 42920 42431 43546
rect 31977 377 32631 1031
rect 33699 -6015 34325 -5389
<< metal4 >>
rect 40086 83905 40742 83906
rect 23903 83904 24557 83905
rect 23903 83252 23904 83904
rect 24556 83252 24557 83904
rect 23903 36393 24557 83252
rect 40086 83251 40087 83905
rect 40741 83251 49583 83905
rect 40086 83250 40742 83251
rect 39924 77721 40580 77722
rect 39924 77067 39925 77721
rect 40579 77067 49095 77721
rect 39924 77066 40580 77067
rect 39762 72179 40418 72180
rect 39762 71525 39763 72179
rect 40417 71525 48933 72179
rect 39762 71524 40418 71525
rect 39682 66315 40338 66316
rect 39682 65661 39683 66315
rect 40337 65661 48771 66315
rect 39682 65660 40338 65661
rect 39762 60213 40418 60214
rect 39762 59559 39763 60213
rect 40417 59559 48285 60213
rect 39762 59558 40418 59559
rect 39762 53707 40418 53708
rect 39762 53053 39763 53707
rect 40417 53053 47879 53707
rect 39762 53052 40418 53053
rect 39518 48165 40174 48166
rect 39518 47511 39519 48165
rect 40173 47511 47473 48165
rect 39518 47510 40174 47511
rect 41804 43546 42432 43547
rect 41804 42920 41805 43546
rect 42431 42920 46973 43546
rect 41804 42919 42432 42920
rect 13117 35739 46905 36393
rect 13117 35413 13771 35739
rect 9910 34759 13771 35413
rect 9910 30162 10564 34759
rect 9904 30161 10570 30162
rect 9904 29497 9905 30161
rect 10569 29497 10570 30161
rect 9904 29496 10570 29497
rect 25150 30119 26004 30286
rect 25150 29465 25251 30119
rect 25905 29465 46905 30119
rect 25150 29286 26004 29465
rect 26380 24079 27036 24080
rect 26380 23425 26381 24079
rect 27035 23425 46905 24079
rect 26380 23424 27036 23425
rect 27514 17961 28170 17962
rect 27514 17307 27515 17961
rect 28169 17307 46825 17961
rect 27514 17306 28170 17307
rect 29056 12239 29712 12240
rect 29056 11585 29057 12239
rect 29711 11585 46825 12239
rect 29056 11584 29712 11585
rect 30318 6341 31226 6508
rect 30318 5687 30435 6341
rect 31089 5687 46581 6341
rect 30318 5550 31226 5687
rect 31884 1031 32792 1180
rect 31884 377 31977 1031
rect 32631 377 46501 1031
rect 31884 222 32792 377
rect 33574 -5389 34450 -5282
rect 33574 -6015 33699 -5389
rect 34325 -6015 46567 -5389
rect 33574 -6138 34450 -6015
use Stage2Pmos  Stage2Pmos_0
timestamp 1670432383
transform 1 0 1960 0 1 53094
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_1
timestamp 1670432383
transform 1 0 2400 0 1 180
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_2
timestamp 1670432383
transform 1 0 2340 0 1 5538
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_3
timestamp 1670432383
transform 1 0 2170 0 1 11354
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_4
timestamp 1670432383
transform 1 0 2094 0 1 17038
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_5
timestamp 1670432383
transform 1 0 2188 0 1 23158
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_6
timestamp 1670432383
transform 1 0 2208 0 1 29240
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_7
timestamp 1670432383
transform 1 0 2112 0 1 35454
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_8
timestamp 1670432383
transform 1 0 2074 0 1 41500
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_9
timestamp 1670432383
transform 1 0 2018 0 1 47392
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_10
timestamp 1670432383
transform 1 0 2036 0 1 82954
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_11
timestamp 1670432383
transform 1 0 1960 0 1 59384
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_12
timestamp 1670432383
transform 1 0 2132 0 1 65448
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_13
timestamp 1670432383
transform 1 0 2132 0 1 71282
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_14
timestamp 1670432383
transform 1 0 2094 0 1 77080
box -2400 -180 7540 5300
use Stage2Pmos  Stage2Pmos_15
timestamp 1670432383
transform 1 0 2520 0 1 -6064
box -2400 -180 7540 5300
<< labels >>
rlabel metal1 -5680 83240 -5054 84024 7 In1
port 0 w
rlabel metal4 40741 83251 49583 83905 3 Y0_I+
port 1 e
rlabel metal1 -5628 77368 -5002 78152 7 In2
port 2 w
rlabel metal4 40579 77067 49095 77721 3 Y0_I-
port 3 e
rlabel metal1 -5588 71568 -4962 72352 7 In3
port 4 w
rlabel metal4 40417 71525 48933 72179 3 Y0_Q+
port 5 e
rlabel metal1 -5588 65742 -4962 66526 7 In4
port 6 w
rlabel metal4 40337 65661 48771 66315 3 Y0_Q-
port 7 e
rlabel metal1 -5746 59680 -5120 60464 7 In5
port 8 w
rlabel metal4 40417 59559 48285 60213 3 Y1_I+
port 9 e
rlabel metal1 -5772 53384 -5146 54168 7 In6
port 10 w
rlabel metal4 40417 53053 47879 53707 3 Y1_I-
port 11 e
rlabel metal1 -5706 47682 -5080 48466 7 In7
port 12 w
rlabel metal4 40173 47511 47473 48165 3 Y1_Q+
port 13 e
rlabel metal1 -5654 41798 -5028 42582 7 In8
port 14 w
rlabel metal4 42431 42920 46973 43546 3 Y1_Q-
port 15 e
rlabel metal1 -5596 35768 -4970 36552 7 In9
port 16 w
rlabel metal4 13117 35739 46905 36393 3 Y2_I+
port 17 e
rlabel metal1 -5510 29526 -4884 30310 7 In10
port 18 w
rlabel metal4 25905 29465 46905 30119 3 Y2_I-
port 19 e
rlabel metal1 -5530 23458 -4904 24242 7 In11
port 20 w
rlabel metal4 27035 23425 46905 24079 3 Y2_Q+
port 21 e
rlabel metal1 -5614 17324 -4988 18108 7 In12
port 22 w
rlabel metal4 28169 17307 46825 17961 3 Y2_Q-
port 23 e
rlabel metal1 -5556 11630 -4930 12414 7 In13
port 24 w
rlabel metal4 29711 11585 46825 12239 3 Y3_I+
port 25 e
rlabel metal1 -5406 5848 -4780 6632 7 In14
port 26 w
rlabel metal4 31089 5687 46581 6341 3 Y3_I-
port 27 e
rlabel metal1 -5322 486 -4696 1270 7 In15
port 28 w
rlabel metal4 32631 377 46501 1031 3 Y3_Q+
port 29 e
rlabel metal1 -4898 -5770 -4272 -4986 7 In16
port 30 w
rlabel metal4 34325 -6015 46567 -5389 3 Y3_Q-
port 31 e
<< end >>
