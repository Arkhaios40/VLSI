magic
tech sky130A
magscale 1 2
timestamp 1670361013
<< nwell >>
rect -558 -1497 558 1497
<< mvpmos >>
rect -300 -1200 300 1200
<< mvpdiff >>
rect -358 1188 -300 1200
rect -358 -1188 -346 1188
rect -312 -1188 -300 1188
rect -358 -1200 -300 -1188
rect 300 1188 358 1200
rect 300 -1188 312 1188
rect 346 -1188 358 1188
rect 300 -1200 358 -1188
<< mvpdiffc >>
rect -346 -1188 -312 1188
rect 312 -1188 346 1188
<< mvnsubdiff >>
rect -492 1419 492 1431
rect -492 1385 -384 1419
rect 384 1385 492 1419
rect -492 1373 492 1385
rect -492 1323 -434 1373
rect -492 -1323 -480 1323
rect -446 -1323 -434 1323
rect 434 1323 492 1373
rect -492 -1373 -434 -1323
rect 434 -1323 446 1323
rect 480 -1323 492 1323
rect 434 -1373 492 -1323
rect -492 -1385 492 -1373
rect -492 -1419 -384 -1385
rect 384 -1419 492 -1385
rect -492 -1431 492 -1419
<< mvnsubdiffcont >>
rect -384 1385 384 1419
rect -480 -1323 -446 1323
rect 446 -1323 480 1323
rect -384 -1419 384 -1385
<< poly >>
rect -300 1281 300 1297
rect -300 1247 -284 1281
rect 284 1247 300 1281
rect -300 1200 300 1247
rect -300 -1247 300 -1200
rect -300 -1281 -284 -1247
rect 284 -1281 300 -1247
rect -300 -1297 300 -1281
<< polycont >>
rect -284 1247 284 1281
rect -284 -1281 284 -1247
<< locali >>
rect -480 1385 -384 1419
rect 384 1385 480 1419
rect -480 1323 -446 1385
rect 446 1323 480 1385
rect -300 1247 -284 1281
rect 284 1247 300 1281
rect -346 1188 -312 1204
rect -346 -1204 -312 -1188
rect 312 1188 346 1204
rect 312 -1204 346 -1188
rect -300 -1281 -284 -1247
rect 284 -1281 300 -1247
rect -480 -1385 -446 -1323
rect 446 -1385 480 -1323
rect -480 -1419 -384 -1385
rect 384 -1419 480 -1385
<< viali >>
rect -284 1247 284 1281
rect -346 -1188 -312 1188
rect 312 -1188 346 1188
rect -284 -1281 284 -1247
<< metal1 >>
rect -296 1281 296 1287
rect -296 1247 -284 1281
rect 284 1247 296 1281
rect -296 1241 296 1247
rect -352 1188 -306 1200
rect -352 -1188 -346 1188
rect -312 -1188 -306 1188
rect -352 -1200 -306 -1188
rect 306 1188 352 1200
rect 306 -1188 312 1188
rect 346 -1188 352 1188
rect 306 -1200 352 -1188
rect -296 -1247 296 -1241
rect -296 -1281 -284 -1247
rect 284 -1281 296 -1247
rect -296 -1287 296 -1281
<< properties >>
string FIXED_BBOX -463 -1402 463 1402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 12 l 3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
