magic
tech sky130A
magscale 1 2
timestamp 1669422754
<< locali >>
rect -1194 13364 268 13366
rect -7176 13348 -5656 13358
rect -7176 12930 -5634 13348
rect -6352 12214 -5634 12930
rect -1202 12918 268 13364
rect -1202 12258 -536 12918
<< viali >>
rect -6352 11496 -5634 12214
rect -1202 11592 -536 12258
<< metal1 >>
rect -1208 12258 -530 12270
rect -6358 12214 -5628 12226
rect -7985 11496 -6352 12214
rect -5634 11496 -5628 12214
rect -1208 11592 -1202 12258
rect -536 11592 -193 12258
rect 473 11592 479 12258
rect -1208 11580 -530 11592
rect -6358 11484 -5628 11496
rect 2521 4690 3111 4696
rect 2521 4094 3111 4100
<< via1 >>
rect -193 11592 473 12258
rect 2521 4100 3111 4690
<< metal2 >>
rect 5652 13250 6308 13259
rect -193 12258 473 12264
rect -193 11093 473 11592
rect 5652 11256 6308 12594
rect 2515 4100 2521 4690
rect 3111 4100 3117 4690
rect 2521 2635 3111 4100
<< via2 >>
rect 5652 12594 6308 13250
<< metal3 >>
rect 5652 13255 6308 13938
rect 5647 13250 6313 13255
rect 5647 12594 5652 13250
rect 6308 12594 6313 13250
rect 5647 12589 6313 12594
use ConnectedNMOSPair  ConnectedNMOSPair_0
timestamp 1669244576
transform 1 0 5644 0 1 4184
box -5846 -84 5646 8110
use CurRefResistor  CurRefResistor_0
timestamp 1669244576
transform 1 0 -9935 0 1 -9501
box 2587 22285 10383 31620
<< labels >>
rlabel metal1 -7985 11496 -6352 12214 7 Vplus
port 0 w
rlabel metal3 5652 13250 6308 13938 1 Ref
port 2 n
rlabel metal2 2521 2635 3111 4100 5 Vneg
port 3 s
<< end >>
