magic
tech sky130A
magscale 1 2
timestamp 1669543272
<< pwell >>
rect -4840 -2540 4080 -2320
<< mvpsubdiff >>
rect -318 -2344 4024 -2332
rect -318 -2360 4028 -2344
rect -340 -2440 4040 -2360
<< locali >>
rect 10440 4720 10800 4780
rect 4120 4560 10800 4720
rect 3340 3440 4280 4380
rect 3340 2920 3620 3440
rect 10440 3260 10800 4560
rect 4120 3100 10800 3260
rect 3340 1980 4280 2920
rect 3340 1460 3620 1980
rect 10440 1800 10800 3100
rect 4120 1640 10800 1800
rect 3340 1360 4280 1460
rect 3122 702 4280 1360
rect 2462 700 4280 702
rect 3340 620 4280 700
rect 3340 520 4020 620
rect 3340 500 3620 520
rect 10440 320 10800 1640
rect 3320 -500 4260 -420
rect 3320 -640 3500 -500
rect 180 -880 3500 -640
rect 4400 -700 9300 -660
rect 4400 -780 4420 -700
rect 4400 -820 9300 -780
rect -4540 -1080 -360 -1040
rect -4540 -1260 -4500 -1080
rect -800 -1260 -360 -1080
rect 180 -1140 240 -880
rect 3220 -980 3500 -880
rect 3220 -1060 4260 -980
rect 3220 -1140 3300 -1060
rect 180 -1220 3300 -1140
rect -4540 -1300 -360 -1260
rect -520 -1344 -360 -1300
rect -478 -1578 -360 -1344
rect -520 -2080 -360 -1578
rect -4520 -2400 -760 -2320
rect -4520 -2520 -4480 -2400
rect -800 -2520 -760 -2400
rect -320 -2344 4020 -2320
rect -320 -2418 4028 -2344
rect -320 -2420 4020 -2418
rect -4520 -2560 -760 -2520
rect 20 -2440 3740 -2420
rect 20 -2540 40 -2440
rect 3720 -2540 3740 -2440
rect 20 -2560 3740 -2540
<< viali >>
rect 10440 4780 10800 5140
rect 2462 702 3122 1360
rect 4420 -780 9300 -700
rect -4500 -1260 -800 -1080
rect 240 -1140 3220 -880
rect -4480 -2520 -800 -2400
rect 40 -2540 3720 -2440
<< metal1 >>
rect 6320 6364 7375 6667
rect 7375 5309 7410 5755
rect 6320 5140 7410 5309
rect 10434 5140 10806 5152
rect 3680 4860 3920 4866
rect 6320 4860 10440 5140
rect 3920 4780 10440 4860
rect 10800 4780 10806 5140
rect 3920 4660 10180 4780
rect 10434 4768 10806 4780
rect 3920 4620 4140 4660
rect 3680 4614 3920 4620
rect 4440 4420 10180 4660
rect 4440 3300 10160 3400
rect -3246 2445 -3240 3195
rect -2490 2445 -2484 3195
rect 10 3165 740 3171
rect -3240 -330 -2490 2445
rect 4440 3060 10880 3300
rect 4440 2960 10160 3060
rect 10 2070 740 2435
rect 1617 2888 2276 2894
rect 2276 2229 3122 2888
rect 1617 2223 2276 2229
rect -40 1452 740 2070
rect -42 642 740 1452
rect 2462 1366 3122 2229
rect 4440 1840 10180 1940
rect 3674 1600 3680 1840
rect 3920 1600 10180 1840
rect 4440 1500 10180 1600
rect 2450 1360 3134 1366
rect 2450 702 2462 1360
rect 3122 702 3134 1360
rect 2450 696 3134 702
rect -3240 -1040 -2460 -330
rect -40 -820 740 642
rect 4380 220 10180 480
rect 3974 -140 3980 220
rect 4340 200 10180 220
rect 10680 200 10880 3060
rect 4340 -120 10660 200
rect 10980 -120 10986 200
rect 4340 -140 9200 -120
rect 4380 -400 9200 -140
rect 4400 -620 9160 -520
rect 4400 -700 9920 -620
rect 4400 -780 4420 -700
rect 9300 -780 9920 -700
rect -40 -880 3380 -820
rect -40 -990 240 -880
rect -4540 -1080 -760 -1040
rect -4540 -1260 -4500 -1080
rect -800 -1260 -760 -1080
rect -176 -1130 -170 -990
rect -30 -1130 240 -990
rect -40 -1140 240 -1130
rect 3220 -1140 3380 -880
rect 4400 -860 9920 -780
rect 4400 -960 9160 -860
rect -40 -1220 3380 -1140
rect -4540 -1560 -760 -1260
rect 0 -1560 3780 -1220
rect 4380 -1340 9200 -1080
rect 4380 -1660 4420 -1340
rect 4740 -1660 9200 -1340
rect 4380 -1700 9200 -1660
rect -4540 -2400 -740 -2180
rect -4540 -2520 -4480 -2400
rect -800 -2520 -740 -2400
rect -4540 -2580 -740 -2520
rect 0 -2440 3760 -2180
rect 0 -2540 40 -2440
rect 3720 -2540 3760 -2440
rect 9580 -2540 9920 -860
rect 0 -2580 9920 -2540
rect -4540 -2760 9920 -2580
rect -650 -4010 -152 -2760
rect 3640 -2780 9920 -2760
rect -650 -4514 -152 -4508
<< via1 >>
rect 6320 5309 7375 6364
rect 3680 4620 3920 4860
rect -3240 2445 -2490 3195
rect 10 2435 740 3165
rect 1617 2229 2276 2888
rect 3680 1600 3920 1840
rect 3980 -140 4340 220
rect 10660 -120 10980 200
rect -170 -1130 -30 -990
rect 4420 -1660 4740 -1340
rect -650 -4508 -152 -4010
<< metal2 >>
rect 6320 6364 7375 8287
rect 6314 5309 6320 6364
rect 7375 5309 7381 6364
rect 3674 4620 3680 4860
rect 3920 4620 3926 4860
rect -3240 3195 -2490 3915
rect 10 3165 740 3925
rect -3240 2439 -2490 2445
rect 4 2435 10 3165
rect 740 2435 746 3165
rect 1617 2888 2276 3993
rect 1611 2229 1617 2888
rect 2276 2229 2282 2888
rect 3680 1840 3920 4620
rect 3680 1594 3920 1600
rect 3980 220 4340 226
rect 3571 -140 3580 220
rect 3940 -140 3980 220
rect 10660 200 10980 206
rect 10980 -120 12280 200
rect 10660 -126 10980 -120
rect 3980 -146 4340 -140
rect -310 -984 -170 -981
rect -310 -990 -30 -984
rect -310 -1136 -30 -1130
rect -310 -1139 -170 -1136
rect 4240 -1310 4780 -1300
rect 4090 -1340 4780 -1310
rect 4090 -1370 4420 -1340
rect 4081 -1700 4090 -1370
rect 4740 -1660 4780 -1340
rect 4420 -1700 4780 -1660
rect -656 -4508 -650 -4010
rect -152 -4508 -146 -4010
rect -650 -5869 -152 -4508
<< via2 >>
rect 3580 -140 3940 220
rect -310 -1130 -170 -990
rect 4090 -1700 4420 -1370
<< metal3 >>
rect 3575 220 3945 225
rect 3074 -140 3080 220
rect 3440 -140 3580 220
rect 3940 -140 3945 220
rect 3575 -145 3945 -140
rect -310 -610 -170 -604
rect -310 -985 -170 -750
rect -315 -990 -165 -985
rect -315 -1130 -310 -990
rect -170 -1130 -165 -990
rect -315 -1135 -165 -1130
rect 4079 -1705 4085 -1365
rect 4410 -1370 4425 -1365
rect 4420 -1700 4425 -1370
rect 4410 -1705 4425 -1700
<< via3 >>
rect 3080 -140 3440 220
rect -310 -750 -170 -610
rect 4085 -1370 4410 -1365
rect 4085 -1700 4090 -1370
rect 4090 -1700 4410 -1370
rect 4085 -1705 4410 -1700
<< metal4 >>
rect -313 540 -166 553
rect -313 -380 240 540
rect 1280 221 3440 540
rect 1280 220 3441 221
rect 1280 -140 3080 220
rect 3440 -140 3441 220
rect 1280 -141 3441 -140
rect 1280 -278 3440 -141
rect 1280 -380 3823 -278
rect -313 -610 -166 -380
rect 2960 -442 3823 -380
rect 3078 -603 3823 -442
rect -313 -750 -310 -610
rect -170 -750 -166 -610
rect -313 -753 -166 -750
rect 3498 -1372 3823 -603
rect 4084 -1365 4411 -1364
rect 4084 -1372 4085 -1365
rect 3498 -1697 4085 -1372
rect 4084 -1705 4085 -1697
rect 4410 -1705 4411 -1365
rect 4084 -1706 4411 -1705
use sky130_fd_pr__cap_mim_m3_1_27X89E  sky130_fd_pr__cap_mim_m3_1_27X89E_0
timestamp 1669447977
transform -1 0 1346 0 -1 80
box -1186 -540 1186 540
use sky130_fd_pr__nfet_g5v0d10v5_2ZQVB2  sky130_fd_pr__nfet_g5v0d10v5_2ZQVB2_0
timestamp 1669452473
transform 0 -1 1847 1 0 -1872
box -528 -2227 528 2447
use sky130_fd_pr__nfet_g5v0d10v5_2ZQVB2  sky130_fd_pr__nfet_g5v0d10v5_2ZQVB2_1
timestamp 1669452473
transform 0 1 -2613 -1 0 -1872
box -528 -2227 528 2447
use sky130_fd_pr__nfet_g5v0d10v5_49CJ6G  sky130_fd_pr__nfet_g5v0d10v5_49CJ6G_0
timestamp 1669438545
transform 0 -1 6767 1 0 -462
box -278 -2727 278 2727
use sky130_fd_pr__nfet_g5v0d10v5_49CJ6G  sky130_fd_pr__nfet_g5v0d10v5_49CJ6G_1
timestamp 1669438545
transform 0 -1 6767 1 0 -1022
box -278 -2727 278 2727
use sky130_fd_pr__pfet_g5v0d10v5_M768YF  sky130_fd_pr__pfet_g5v0d10v5_M768YF_0
timestamp 1669447977
transform 0 -1 7322 1 0 3938
box -758 -3262 758 3262
use sky130_fd_pr__pfet_g5v0d10v5_M768YF  sky130_fd_pr__pfet_g5v0d10v5_M768YF_1
timestamp 1669447977
transform 0 -1 7322 1 0 2478
box -758 -3262 758 3262
use sky130_fd_pr__pfet_g5v0d10v5_M768YF  sky130_fd_pr__pfet_g5v0d10v5_M768YF_2
timestamp 1669447977
transform 0 -1 7322 1 0 1018
box -758 -3262 758 3262
<< labels >>
rlabel metal2 6820 7900 6820 7900 1 VPlus
port 0 n
rlabel metal2 -2900 3700 -2900 3700 1 Gain_L_Pin
port 1 n
rlabel metal2 340 3740 340 3740 1 Gain_R_Pin
port 2 n
rlabel metal1 9500 -760 9500 -760 1 1
rlabel metal2 1617 2888 2276 3993 1 GateRef
port 3 n
rlabel metal2 10980 -120 12280 200 3 Out
port 4 e
rlabel metal2 -650 -5869 -152 -4508 5 Gain_Vs
port 5 s
<< end >>
