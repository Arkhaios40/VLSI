** sch_path: /home/arkhaios/Project/xschem/PrimalStructures/Level2/CurrentRef.sch
**.subckt CurrentRef Vplus Body Ref Vneg
*.iopin Vplus
*.iopin Body
*.iopin Ref
*.iopin Vneg
x6 Vplus Body net1 CurRefResistor
x1 Ref net1 Vneg ConnectedNMOSPair
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  PrimalStructures/CurRefResistor.sym # of pins=3
** sym_path: /home/arkhaios/Project/xschem/PrimalStructures/CurRefResistor.sym
** sch_path: /home/arkhaios/Project/xschem/PrimalStructures/CurRefResistor.sch
.subckt CurRefResistor Pin1 Body Pin2
*.iopin Pin1
*.iopin Pin2
*.iopin Body
XR1 Pin2 Pin1 Body sky130_fd_pr__res_xhigh_po_1p41 L=40 mult=1 m=1
.ends


* expanding   symbol:  PrimalStructures/Level2/ConnectedNMOSPair.sym # of pins=3
** sym_path: /home/arkhaios/Project/xschem/PrimalStructures/Level2/ConnectedNMOSPair.sym
** sch_path: /home/arkhaios/Project/xschem/PrimalStructures/Level2/ConnectedNMOSPair.sch
.subckt ConnectedNMOSPair R_Pin L_Pin Vs
*.iopin L_Pin
*.iopin R_Pin
*.iopin Vs
x1 L_Pin L_Pin Vs Vs NMOSPair
x2 R_Pin L_Pin Vs Vs NMOSPair
.ends


* expanding   symbol:  PrimalStructures/NMOSPair.sym # of pins=4
** sym_path: /home/arkhaios/Project/xschem/PrimalStructures/NMOSPair.sym
** sch_path: /home/arkhaios/Project/xschem/PrimalStructures/NMOSPair.sch
.subckt NMOSPair Vd Vn Vnbody Vs
*.iopin Vd
*.iopin Vn
*.iopin Vnbody
*.iopin Vs
XM1 Vd Vn net1 Vnbody sky130_fd_pr__nfet_g5v0d10v5 L=2 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vd Vn net1 Vnbody sky130_fd_pr__nfet_g5v0d10v5 L=2 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vd Vn net1 Vnbody sky130_fd_pr__nfet_g5v0d10v5 L=2 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 Vd Vn net1 Vnbody sky130_fd_pr__nfet_g5v0d10v5 L=2 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vd Vn net1 Vnbody sky130_fd_pr__nfet_g5v0d10v5 L=2 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net1 Vn Vs Vnbody sky130_fd_pr__nfet_g5v0d10v5 L=5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
