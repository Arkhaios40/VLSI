magic
tech sky130A
magscale 1 2
timestamp 1668639803
<< nwell >>
rect -758 -3297 758 3297
<< mvpmos >>
rect -500 -3000 500 3000
<< mvpdiff >>
rect -558 2988 -500 3000
rect -558 -2988 -546 2988
rect -512 -2988 -500 2988
rect -558 -3000 -500 -2988
rect 500 2988 558 3000
rect 500 -2988 512 2988
rect 546 -2988 558 2988
rect 500 -3000 558 -2988
<< mvpdiffc >>
rect -546 -2988 -512 2988
rect 512 -2988 546 2988
<< mvnsubdiff >>
rect -692 3173 692 3231
rect -692 3123 -634 3173
rect -692 -3123 -680 3123
rect -646 -3123 -634 3123
rect 634 3123 692 3173
rect -692 -3173 -634 -3123
rect 634 -3123 646 3123
rect 680 -3123 692 3123
rect 634 -3173 692 -3123
rect -692 -3231 692 -3173
<< mvnsubdiffcont >>
rect -680 -3123 -646 3123
rect 646 -3123 680 3123
<< poly >>
rect -500 3000 500 3097
rect -500 -3047 500 -3000
rect -500 -3081 -484 -3047
rect 484 -3081 500 -3047
rect -500 -3097 500 -3081
<< polycont >>
rect -484 -3081 484 -3047
<< locali >>
rect -680 3123 -646 3157
rect 646 3123 680 3157
rect -546 2988 -512 3004
rect -546 -3004 -512 -2988
rect 512 2988 546 3004
rect 512 -3005 546 -2988
rect -500 -3081 -484 -3047
rect 484 -3081 500 -3047
rect -680 -3145 -646 -3123
rect 646 -3145 680 -3123
<< viali >>
rect -546 -2988 -512 2988
rect 512 -2988 546 2988
rect -484 -3081 484 -3047
<< metal1 >>
rect -552 2988 -506 3000
rect -552 -2988 -546 2988
rect -512 -2988 -506 2988
rect -552 -3000 -506 -2988
rect 506 2988 552 3000
rect 506 -2988 512 2988
rect 546 -2988 552 2988
rect 506 -3000 552 -2988
rect -496 -3047 496 -3041
rect -496 -3081 -484 -3047
rect 484 -3081 496 -3047
rect -496 -3087 496 -3081
<< properties >>
string FIXED_BBOX -663 -3202 663 3202
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 30.0 l 5.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
