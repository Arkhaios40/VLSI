magic
tech sky130A
magscale 1 2
timestamp 1670358787
<< checkpaint >>
rect -1260 -660 7271 6111
rect -1260 -2346 1460 -660
rect -1260 -7660 39193 -2346
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
use NmosStage1  NmosStage1_0
timestamp 1670353092
transform 1 0 65 0 1 1400
box 0 -800 5419 1994
use NmosStage1  x1
timestamp 1670353092
transform 1 0 0 0 1 -5600
box 0 -800 5419 1994
use NmosStage1  x3
timestamp 1670353092
transform 1 0 5419 0 1 -5600
box 0 -800 5419 1994
use NmosStage1  x4
timestamp 1670353092
transform 1 0 10838 0 1 -5600
box 0 -800 5419 1994
use NmosStage1  x5
timestamp 1670353092
transform 1 0 16257 0 1 -5600
box 0 -800 5419 1994
use NmosStage1  x6
timestamp 1670353092
transform 1 0 21676 0 1 -5600
box 0 -800 5419 1994
use NmosStage1  x7
timestamp 1670353092
transform 1 0 27095 0 1 -5600
box 0 -800 5419 1994
use NmosStage1  x8
timestamp 1670353092
transform 1 0 32514 0 1 -5600
box 0 -800 5419 1994
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 IN_X0_i+
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Out1
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 IN_X0_i-
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Out2
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 IN_X0_q+
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Out3
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 IN_X0_q-
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 Out4
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 IN_X2_i+
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 Out5
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 IN_X2_i-
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 {}
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 Out6
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 IN_X2_q+
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 Out7
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 IN_X2_q-
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 Out8
port 16 nsew
<< end >>
